module linear_DW01_add_21 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [7:1] carry;

  FADDX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FADDX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FADDX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FADDX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(n1), .CO(carry[3]), .S(SUM[2]) );
  INVX0 U1 ( .INP(carry[6]), .ZN(n4) );
  NAND2X1 U2 ( .IN1(n3), .IN2(n4), .QN(carry[7]) );
  INVX0 U3 ( .INP(B[6]), .ZN(n3) );
  AND2X1 U4 ( .IN1(B[1]), .IN2(n2), .Q(n1) );
  AND2X1 U5 ( .IN1(B[0]), .IN2(CI), .Q(n2) );
  XOR2X1 U6 ( .IN1(n4), .IN2(B[6]), .Q(SUM[6]) );
  XOR2X1 U7 ( .IN1(B[7]), .IN2(carry[7]), .Q(SUM[7]) );
  XOR2X1 U8 ( .IN1(B[1]), .IN2(n2), .Q(SUM[1]) );
  XOR2X1 U9 ( .IN1(B[0]), .IN2(CI), .Q(SUM[0]) );
endmodule


module linear_DW01_add_23 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [7:1] carry;

  FADDX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FADDX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FADDX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FADDX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(n1), .CO(carry[3]), .S(SUM[2]) );
  INVX0 U1 ( .INP(carry[6]), .ZN(n4) );
  NAND2X1 U2 ( .IN1(n3), .IN2(n4), .QN(carry[7]) );
  INVX0 U3 ( .INP(B[6]), .ZN(n3) );
  AND2X1 U4 ( .IN1(B[1]), .IN2(n2), .Q(n1) );
  AND2X1 U5 ( .IN1(B[0]), .IN2(CI), .Q(n2) );
  XOR2X1 U6 ( .IN1(n4), .IN2(B[6]), .Q(SUM[6]) );
  XOR2X1 U7 ( .IN1(B[7]), .IN2(carry[7]), .Q(SUM[7]) );
  XOR2X1 U8 ( .IN1(B[1]), .IN2(n2), .Q(SUM[1]) );
  XOR2X1 U9 ( .IN1(B[0]), .IN2(CI), .Q(SUM[0]) );
endmodule


module linear_DW01_add_25 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [7:1] carry;

  FADDX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FADDX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FADDX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FADDX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(n1), .CO(carry[3]), .S(SUM[2]) );
  INVX0 U1 ( .INP(carry[6]), .ZN(n4) );
  NAND2X1 U2 ( .IN1(n3), .IN2(n4), .QN(carry[7]) );
  INVX0 U3 ( .INP(B[6]), .ZN(n3) );
  AND2X1 U4 ( .IN1(B[1]), .IN2(n2), .Q(n1) );
  AND2X1 U5 ( .IN1(B[0]), .IN2(CI), .Q(n2) );
  XOR2X1 U6 ( .IN1(n4), .IN2(B[6]), .Q(SUM[6]) );
  XOR2X1 U7 ( .IN1(B[7]), .IN2(carry[7]), .Q(SUM[7]) );
  XOR2X1 U8 ( .IN1(B[1]), .IN2(n2), .Q(SUM[1]) );
  XOR2X1 U9 ( .IN1(B[0]), .IN2(CI), .Q(SUM[0]) );
endmodule


module linear_DW01_add_27 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [7:1] carry;

  FADDX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FADDX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FADDX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FADDX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(n1), .CO(carry[3]), .S(SUM[2]) );
  INVX0 U1 ( .INP(carry[6]), .ZN(n4) );
  NAND2X1 U2 ( .IN1(n3), .IN2(n4), .QN(carry[7]) );
  INVX0 U3 ( .INP(B[6]), .ZN(n3) );
  AND2X1 U4 ( .IN1(B[1]), .IN2(n2), .Q(n1) );
  AND2X1 U5 ( .IN1(B[0]), .IN2(CI), .Q(n2) );
  XOR2X1 U6 ( .IN1(n4), .IN2(B[6]), .Q(SUM[6]) );
  XOR2X1 U7 ( .IN1(B[7]), .IN2(carry[7]), .Q(SUM[7]) );
  XOR2X1 U8 ( .IN1(B[1]), .IN2(n2), .Q(SUM[1]) );
  XOR2X1 U9 ( .IN1(B[0]), .IN2(CI), .Q(SUM[0]) );
endmodule


module linear_DW01_add_29 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [7:1] carry;

  FADDX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FADDX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FADDX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FADDX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(n1), .CO(carry[3]), .S(SUM[2]) );
  INVX0 U1 ( .INP(carry[6]), .ZN(n4) );
  NAND2X1 U2 ( .IN1(n3), .IN2(n4), .QN(carry[7]) );
  INVX0 U3 ( .INP(B[6]), .ZN(n3) );
  AND2X1 U4 ( .IN1(B[1]), .IN2(n2), .Q(n1) );
  AND2X1 U5 ( .IN1(B[0]), .IN2(CI), .Q(n2) );
  XOR2X1 U6 ( .IN1(n4), .IN2(B[6]), .Q(SUM[6]) );
  XOR2X1 U7 ( .IN1(B[7]), .IN2(carry[7]), .Q(SUM[7]) );
  XOR2X1 U8 ( .IN1(B[1]), .IN2(n2), .Q(SUM[1]) );
  XOR2X1 U9 ( .IN1(B[0]), .IN2(CI), .Q(SUM[0]) );
endmodule


module linear_DW01_add_31 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [7:1] carry;

  FADDX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FADDX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FADDX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FADDX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(n1), .CO(carry[3]), .S(SUM[2]) );
  INVX0 U1 ( .INP(carry[6]), .ZN(n4) );
  NAND2X1 U2 ( .IN1(n3), .IN2(n4), .QN(carry[7]) );
  INVX0 U3 ( .INP(B[6]), .ZN(n3) );
  AND2X1 U4 ( .IN1(B[1]), .IN2(n2), .Q(n1) );
  AND2X1 U5 ( .IN1(B[0]), .IN2(CI), .Q(n2) );
  XOR2X1 U6 ( .IN1(n4), .IN2(B[6]), .Q(SUM[6]) );
  XOR2X1 U7 ( .IN1(B[7]), .IN2(carry[7]), .Q(SUM[7]) );
  XOR2X1 U8 ( .IN1(B[1]), .IN2(n2), .Q(SUM[1]) );
  XOR2X1 U9 ( .IN1(B[0]), .IN2(CI), .Q(SUM[0]) );
endmodule


module linear_DW01_add_33 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [7:1] carry;

  FADDX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FADDX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FADDX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FADDX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(n1), .CO(carry[3]), .S(SUM[2]) );
  INVX0 U1 ( .INP(carry[6]), .ZN(n4) );
  NAND2X1 U2 ( .IN1(n3), .IN2(n4), .QN(carry[7]) );
  INVX0 U3 ( .INP(B[6]), .ZN(n3) );
  AND2X1 U4 ( .IN1(B[1]), .IN2(n2), .Q(n1) );
  AND2X1 U5 ( .IN1(B[0]), .IN2(CI), .Q(n2) );
  XOR2X1 U6 ( .IN1(n4), .IN2(B[6]), .Q(SUM[6]) );
  XOR2X1 U7 ( .IN1(B[7]), .IN2(carry[7]), .Q(SUM[7]) );
  XOR2X1 U8 ( .IN1(B[1]), .IN2(n2), .Q(SUM[1]) );
  XOR2X1 U9 ( .IN1(B[0]), .IN2(CI), .Q(SUM[0]) );
endmodule


module linear_DW01_add_35 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [7:1] carry;

  FADDX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FADDX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FADDX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FADDX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(n1), .CO(carry[3]), .S(SUM[2]) );
  INVX0 U1 ( .INP(carry[6]), .ZN(n4) );
  NAND2X1 U2 ( .IN1(n3), .IN2(n4), .QN(carry[7]) );
  INVX0 U3 ( .INP(B[6]), .ZN(n3) );
  AND2X1 U4 ( .IN1(B[1]), .IN2(n2), .Q(n1) );
  AND2X1 U5 ( .IN1(B[0]), .IN2(CI), .Q(n2) );
  XOR2X1 U6 ( .IN1(n4), .IN2(B[6]), .Q(SUM[6]) );
  XOR2X1 U7 ( .IN1(B[7]), .IN2(carry[7]), .Q(SUM[7]) );
  XOR2X1 U8 ( .IN1(B[1]), .IN2(n2), .Q(SUM[1]) );
  XOR2X1 U9 ( .IN1(B[0]), .IN2(CI), .Q(SUM[0]) );
endmodule


module linear_DW01_add_37 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [7:1] carry;

  FADDX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FADDX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FADDX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FADDX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(n1), .CO(carry[3]), .S(SUM[2]) );
  INVX0 U1 ( .INP(carry[6]), .ZN(n4) );
  NAND2X1 U2 ( .IN1(n3), .IN2(n4), .QN(carry[7]) );
  INVX0 U3 ( .INP(B[6]), .ZN(n3) );
  AND2X1 U4 ( .IN1(B[1]), .IN2(n2), .Q(n1) );
  AND2X1 U5 ( .IN1(B[0]), .IN2(CI), .Q(n2) );
  XOR2X1 U6 ( .IN1(n4), .IN2(B[6]), .Q(SUM[6]) );
  XOR2X1 U7 ( .IN1(B[7]), .IN2(carry[7]), .Q(SUM[7]) );
  XOR2X1 U8 ( .IN1(B[1]), .IN2(n2), .Q(SUM[1]) );
  XOR2X1 U9 ( .IN1(B[0]), .IN2(CI), .Q(SUM[0]) );
endmodule


module linear_DW01_add_39 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [7:1] carry;

  FADDX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FADDX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FADDX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FADDX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(n1), .CO(carry[3]), .S(SUM[2]) );
  INVX0 U1 ( .INP(carry[6]), .ZN(n4) );
  NAND2X1 U2 ( .IN1(n3), .IN2(n4), .QN(carry[7]) );
  INVX0 U3 ( .INP(B[6]), .ZN(n3) );
  AND2X1 U4 ( .IN1(B[1]), .IN2(n2), .Q(n1) );
  AND2X1 U5 ( .IN1(B[0]), .IN2(CI), .Q(n2) );
  XOR2X1 U6 ( .IN1(n4), .IN2(B[6]), .Q(SUM[6]) );
  XOR2X1 U7 ( .IN1(B[7]), .IN2(carry[7]), .Q(SUM[7]) );
  XOR2X1 U8 ( .IN1(B[1]), .IN2(n2), .Q(SUM[1]) );
  XOR2X1 U9 ( .IN1(B[0]), .IN2(CI), .Q(SUM[0]) );
endmodule


module linear_DW_mult_uns_0 ( a, b, product );
  input [4:0] a;
  input [4:0] b;
  output [9:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n89, n90, n91,
         n92, n93, n94, n95, n96;
  assign n33 = b[3];
  assign n34 = b[2];
  assign n35 = b[1];
  assign n36 = b[0];
  assign n37 = a[3];
  assign n42 = a[2];
  assign n47 = a[1];
  assign n52 = a[0];

  FADDX1 U4 ( .A(n11), .B(n10), .CI(n3), .CO(n2), .S(product[7]) );
  FADDX1 U5 ( .A(n12), .B(n15), .CI(n4), .CO(n3), .S(product[6]) );
  FADDX1 U6 ( .A(n16), .B(n21), .CI(n5), .CO(n4), .S(product[5]) );
  FADDX1 U7 ( .A(n22), .B(n27), .CI(n6), .CO(n5), .S(product[4]) );
  FADDX1 U8 ( .A(n28), .B(n31), .CI(n7), .CO(n6), .S(product[3]) );
  FADDX1 U9 ( .A(n32), .B(n46), .CI(n8), .CO(n7), .S(product[2]) );
  HADDX1 U10 ( .A0(n51), .B0(n55), .C1(n8), .SO(product[1]) );
  FADDX1 U11 ( .A(n33), .B(n37), .CI(n13), .CO(n9), .S(n10) );
  FADDX1 U12 ( .A(n14), .B(n19), .CI(n17), .CO(n11), .S(n12) );
  FADDX1 U13 ( .A(n34), .B(n42), .CI(n38), .CO(n13), .S(n14) );
  FADDX1 U14 ( .A(n23), .B(n25), .CI(n18), .CO(n15), .S(n16) );
  FADDX1 U15 ( .A(n39), .B(n43), .CI(n20), .CO(n17), .S(n18) );
  HADDX1 U16 ( .A0(n47), .B0(n35), .C1(n19), .SO(n20) );
  FADDX1 U17 ( .A(n29), .B(n26), .CI(n24), .CO(n21), .S(n22) );
  FADDX1 U18 ( .A(n40), .B(n48), .CI(n44), .CO(n23), .S(n24) );
  HADDX1 U19 ( .A0(n36), .B0(n52), .C1(n25), .SO(n26) );
  FADDX1 U20 ( .A(n49), .B(n53), .CI(n30), .CO(n27), .S(n28) );
  HADDX1 U21 ( .A0(n45), .B0(n41), .C1(n29), .SO(n30) );
  HADDX1 U22 ( .A0(n54), .B0(n50), .C1(n31), .SO(n32) );
  INVX0 U58 ( .INP(n34), .ZN(n90) );
  INVX0 U59 ( .INP(n42), .ZN(n94) );
  INVX0 U60 ( .INP(n37), .ZN(n93) );
  INVX0 U61 ( .INP(n52), .ZN(n96) );
  INVX0 U62 ( .INP(n47), .ZN(n95) );
  INVX0 U63 ( .INP(n33), .ZN(n89) );
  INVX0 U64 ( .INP(n35), .ZN(n91) );
  INVX0 U65 ( .INP(n36), .ZN(n92) );
  OR2X1 U66 ( .IN1(n2), .IN2(n9), .Q(product[9]) );
  XNOR2X1 U67 ( .IN1(n2), .IN2(n9), .Q(product[8]) );
  NOR2X0 U68 ( .IN1(n96), .IN2(n92), .QN(product[0]) );
  NOR2X0 U69 ( .IN1(n96), .IN2(n91), .QN(n55) );
  NOR2X0 U70 ( .IN1(n96), .IN2(n90), .QN(n54) );
  NOR2X0 U71 ( .IN1(n96), .IN2(n89), .QN(n53) );
  NOR2X0 U72 ( .IN1(n92), .IN2(n95), .QN(n51) );
  NOR2X0 U73 ( .IN1(n91), .IN2(n95), .QN(n50) );
  NOR2X0 U74 ( .IN1(n90), .IN2(n95), .QN(n49) );
  NOR2X0 U75 ( .IN1(n89), .IN2(n95), .QN(n48) );
  NOR2X0 U76 ( .IN1(n92), .IN2(n94), .QN(n46) );
  NOR2X0 U77 ( .IN1(n91), .IN2(n94), .QN(n45) );
  NOR2X0 U78 ( .IN1(n90), .IN2(n94), .QN(n44) );
  NOR2X0 U79 ( .IN1(n89), .IN2(n94), .QN(n43) );
  NOR2X0 U80 ( .IN1(n92), .IN2(n93), .QN(n41) );
  NOR2X0 U81 ( .IN1(n91), .IN2(n93), .QN(n40) );
  NOR2X0 U82 ( .IN1(n90), .IN2(n93), .QN(n39) );
  NOR2X0 U83 ( .IN1(n89), .IN2(n93), .QN(n38) );
endmodule


module linear_DW_mult_uns_1 ( a, b, product );
  input [4:0] a;
  input [4:0] b;
  output [9:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n89, n90, n91,
         n92, n93, n94, n95, n96;
  assign n33 = b[3];
  assign n34 = b[2];
  assign n35 = b[1];
  assign n36 = b[0];
  assign n37 = a[3];
  assign n42 = a[2];
  assign n47 = a[1];
  assign n52 = a[0];

  FADDX1 U4 ( .A(n11), .B(n10), .CI(n3), .CO(n2), .S(product[7]) );
  FADDX1 U5 ( .A(n12), .B(n15), .CI(n4), .CO(n3), .S(product[6]) );
  FADDX1 U6 ( .A(n16), .B(n21), .CI(n5), .CO(n4), .S(product[5]) );
  FADDX1 U7 ( .A(n22), .B(n27), .CI(n6), .CO(n5), .S(product[4]) );
  FADDX1 U8 ( .A(n28), .B(n31), .CI(n7), .CO(n6), .S(product[3]) );
  FADDX1 U9 ( .A(n32), .B(n46), .CI(n8), .CO(n7), .S(product[2]) );
  HADDX1 U10 ( .A0(n51), .B0(n55), .C1(n8), .SO(product[1]) );
  FADDX1 U11 ( .A(n33), .B(n37), .CI(n13), .CO(n9), .S(n10) );
  FADDX1 U12 ( .A(n14), .B(n19), .CI(n17), .CO(n11), .S(n12) );
  FADDX1 U13 ( .A(n34), .B(n42), .CI(n38), .CO(n13), .S(n14) );
  FADDX1 U14 ( .A(n23), .B(n25), .CI(n18), .CO(n15), .S(n16) );
  FADDX1 U15 ( .A(n39), .B(n43), .CI(n20), .CO(n17), .S(n18) );
  HADDX1 U16 ( .A0(n47), .B0(n35), .C1(n19), .SO(n20) );
  FADDX1 U17 ( .A(n29), .B(n26), .CI(n24), .CO(n21), .S(n22) );
  FADDX1 U18 ( .A(n40), .B(n48), .CI(n44), .CO(n23), .S(n24) );
  HADDX1 U19 ( .A0(n36), .B0(n52), .C1(n25), .SO(n26) );
  FADDX1 U20 ( .A(n49), .B(n53), .CI(n30), .CO(n27), .S(n28) );
  HADDX1 U21 ( .A0(n45), .B0(n41), .C1(n29), .SO(n30) );
  HADDX1 U22 ( .A0(n54), .B0(n50), .C1(n31), .SO(n32) );
  INVX0 U58 ( .INP(n34), .ZN(n90) );
  INVX0 U59 ( .INP(n42), .ZN(n94) );
  INVX0 U60 ( .INP(n37), .ZN(n93) );
  INVX0 U61 ( .INP(n52), .ZN(n96) );
  INVX0 U62 ( .INP(n47), .ZN(n95) );
  INVX0 U63 ( .INP(n33), .ZN(n89) );
  INVX0 U64 ( .INP(n35), .ZN(n91) );
  INVX0 U65 ( .INP(n36), .ZN(n92) );
  OR2X1 U66 ( .IN1(n2), .IN2(n9), .Q(product[9]) );
  XNOR2X1 U67 ( .IN1(n2), .IN2(n9), .Q(product[8]) );
  NOR2X0 U68 ( .IN1(n96), .IN2(n92), .QN(product[0]) );
  NOR2X0 U69 ( .IN1(n96), .IN2(n91), .QN(n55) );
  NOR2X0 U70 ( .IN1(n96), .IN2(n90), .QN(n54) );
  NOR2X0 U71 ( .IN1(n96), .IN2(n89), .QN(n53) );
  NOR2X0 U72 ( .IN1(n92), .IN2(n95), .QN(n51) );
  NOR2X0 U73 ( .IN1(n91), .IN2(n95), .QN(n50) );
  NOR2X0 U74 ( .IN1(n90), .IN2(n95), .QN(n49) );
  NOR2X0 U75 ( .IN1(n89), .IN2(n95), .QN(n48) );
  NOR2X0 U76 ( .IN1(n92), .IN2(n94), .QN(n46) );
  NOR2X0 U77 ( .IN1(n91), .IN2(n94), .QN(n45) );
  NOR2X0 U78 ( .IN1(n90), .IN2(n94), .QN(n44) );
  NOR2X0 U79 ( .IN1(n89), .IN2(n94), .QN(n43) );
  NOR2X0 U80 ( .IN1(n92), .IN2(n93), .QN(n41) );
  NOR2X0 U81 ( .IN1(n91), .IN2(n93), .QN(n40) );
  NOR2X0 U82 ( .IN1(n90), .IN2(n93), .QN(n39) );
  NOR2X0 U83 ( .IN1(n89), .IN2(n93), .QN(n38) );
endmodule


module linear_DW_mult_uns_2 ( a, b, product );
  input [4:0] a;
  input [4:0] b;
  output [9:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n89, n90, n91,
         n92, n93, n94, n95, n96;
  assign n33 = b[3];
  assign n34 = b[2];
  assign n35 = b[1];
  assign n36 = b[0];
  assign n37 = a[3];
  assign n42 = a[2];
  assign n47 = a[1];
  assign n52 = a[0];

  FADDX1 U4 ( .A(n11), .B(n10), .CI(n3), .CO(n2), .S(product[7]) );
  FADDX1 U5 ( .A(n12), .B(n15), .CI(n4), .CO(n3), .S(product[6]) );
  FADDX1 U6 ( .A(n16), .B(n21), .CI(n5), .CO(n4), .S(product[5]) );
  FADDX1 U7 ( .A(n22), .B(n27), .CI(n6), .CO(n5), .S(product[4]) );
  FADDX1 U8 ( .A(n28), .B(n31), .CI(n7), .CO(n6), .S(product[3]) );
  FADDX1 U9 ( .A(n32), .B(n46), .CI(n8), .CO(n7), .S(product[2]) );
  HADDX1 U10 ( .A0(n51), .B0(n55), .C1(n8), .SO(product[1]) );
  FADDX1 U11 ( .A(n33), .B(n37), .CI(n13), .CO(n9), .S(n10) );
  FADDX1 U12 ( .A(n14), .B(n19), .CI(n17), .CO(n11), .S(n12) );
  FADDX1 U13 ( .A(n34), .B(n42), .CI(n38), .CO(n13), .S(n14) );
  FADDX1 U14 ( .A(n23), .B(n25), .CI(n18), .CO(n15), .S(n16) );
  FADDX1 U15 ( .A(n39), .B(n43), .CI(n20), .CO(n17), .S(n18) );
  HADDX1 U16 ( .A0(n47), .B0(n35), .C1(n19), .SO(n20) );
  FADDX1 U17 ( .A(n29), .B(n26), .CI(n24), .CO(n21), .S(n22) );
  FADDX1 U18 ( .A(n40), .B(n48), .CI(n44), .CO(n23), .S(n24) );
  HADDX1 U19 ( .A0(n36), .B0(n52), .C1(n25), .SO(n26) );
  FADDX1 U20 ( .A(n49), .B(n53), .CI(n30), .CO(n27), .S(n28) );
  HADDX1 U21 ( .A0(n45), .B0(n41), .C1(n29), .SO(n30) );
  HADDX1 U22 ( .A0(n54), .B0(n50), .C1(n31), .SO(n32) );
  INVX0 U58 ( .INP(n34), .ZN(n90) );
  INVX0 U59 ( .INP(n42), .ZN(n94) );
  INVX0 U60 ( .INP(n37), .ZN(n93) );
  INVX0 U61 ( .INP(n52), .ZN(n96) );
  INVX0 U62 ( .INP(n47), .ZN(n95) );
  INVX0 U63 ( .INP(n33), .ZN(n89) );
  INVX0 U64 ( .INP(n35), .ZN(n91) );
  INVX0 U65 ( .INP(n36), .ZN(n92) );
  OR2X1 U66 ( .IN1(n2), .IN2(n9), .Q(product[9]) );
  XNOR2X1 U67 ( .IN1(n2), .IN2(n9), .Q(product[8]) );
  NOR2X0 U68 ( .IN1(n96), .IN2(n92), .QN(product[0]) );
  NOR2X0 U69 ( .IN1(n96), .IN2(n91), .QN(n55) );
  NOR2X0 U70 ( .IN1(n96), .IN2(n90), .QN(n54) );
  NOR2X0 U71 ( .IN1(n96), .IN2(n89), .QN(n53) );
  NOR2X0 U72 ( .IN1(n92), .IN2(n95), .QN(n51) );
  NOR2X0 U73 ( .IN1(n91), .IN2(n95), .QN(n50) );
  NOR2X0 U74 ( .IN1(n90), .IN2(n95), .QN(n49) );
  NOR2X0 U75 ( .IN1(n89), .IN2(n95), .QN(n48) );
  NOR2X0 U76 ( .IN1(n92), .IN2(n94), .QN(n46) );
  NOR2X0 U77 ( .IN1(n91), .IN2(n94), .QN(n45) );
  NOR2X0 U78 ( .IN1(n90), .IN2(n94), .QN(n44) );
  NOR2X0 U79 ( .IN1(n89), .IN2(n94), .QN(n43) );
  NOR2X0 U80 ( .IN1(n92), .IN2(n93), .QN(n41) );
  NOR2X0 U81 ( .IN1(n91), .IN2(n93), .QN(n40) );
  NOR2X0 U82 ( .IN1(n90), .IN2(n93), .QN(n39) );
  NOR2X0 U83 ( .IN1(n89), .IN2(n93), .QN(n38) );
endmodule


module linear_DW_mult_uns_3 ( a, b, product );
  input [4:0] a;
  input [4:0] b;
  output [9:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n89, n90, n91,
         n92, n93, n94, n95, n96;
  assign n33 = b[3];
  assign n34 = b[2];
  assign n35 = b[1];
  assign n36 = b[0];
  assign n37 = a[3];
  assign n42 = a[2];
  assign n47 = a[1];
  assign n52 = a[0];

  FADDX1 U4 ( .A(n11), .B(n10), .CI(n3), .CO(n2), .S(product[7]) );
  FADDX1 U5 ( .A(n12), .B(n15), .CI(n4), .CO(n3), .S(product[6]) );
  FADDX1 U6 ( .A(n16), .B(n21), .CI(n5), .CO(n4), .S(product[5]) );
  FADDX1 U7 ( .A(n22), .B(n27), .CI(n6), .CO(n5), .S(product[4]) );
  FADDX1 U8 ( .A(n28), .B(n31), .CI(n7), .CO(n6), .S(product[3]) );
  FADDX1 U9 ( .A(n32), .B(n46), .CI(n8), .CO(n7), .S(product[2]) );
  HADDX1 U10 ( .A0(n51), .B0(n55), .C1(n8), .SO(product[1]) );
  FADDX1 U11 ( .A(n33), .B(n37), .CI(n13), .CO(n9), .S(n10) );
  FADDX1 U12 ( .A(n14), .B(n19), .CI(n17), .CO(n11), .S(n12) );
  FADDX1 U13 ( .A(n34), .B(n42), .CI(n38), .CO(n13), .S(n14) );
  FADDX1 U14 ( .A(n23), .B(n25), .CI(n18), .CO(n15), .S(n16) );
  FADDX1 U15 ( .A(n39), .B(n43), .CI(n20), .CO(n17), .S(n18) );
  HADDX1 U16 ( .A0(n47), .B0(n35), .C1(n19), .SO(n20) );
  FADDX1 U17 ( .A(n29), .B(n26), .CI(n24), .CO(n21), .S(n22) );
  FADDX1 U18 ( .A(n40), .B(n48), .CI(n44), .CO(n23), .S(n24) );
  HADDX1 U19 ( .A0(n36), .B0(n52), .C1(n25), .SO(n26) );
  FADDX1 U20 ( .A(n49), .B(n53), .CI(n30), .CO(n27), .S(n28) );
  HADDX1 U21 ( .A0(n45), .B0(n41), .C1(n29), .SO(n30) );
  HADDX1 U22 ( .A0(n54), .B0(n50), .C1(n31), .SO(n32) );
  INVX0 U58 ( .INP(n34), .ZN(n90) );
  INVX0 U59 ( .INP(n42), .ZN(n94) );
  INVX0 U60 ( .INP(n37), .ZN(n93) );
  INVX0 U61 ( .INP(n52), .ZN(n96) );
  INVX0 U62 ( .INP(n47), .ZN(n95) );
  INVX0 U63 ( .INP(n33), .ZN(n89) );
  INVX0 U64 ( .INP(n35), .ZN(n91) );
  INVX0 U65 ( .INP(n36), .ZN(n92) );
  OR2X1 U66 ( .IN1(n2), .IN2(n9), .Q(product[9]) );
  XNOR2X1 U67 ( .IN1(n2), .IN2(n9), .Q(product[8]) );
  NOR2X0 U68 ( .IN1(n96), .IN2(n92), .QN(product[0]) );
  NOR2X0 U69 ( .IN1(n96), .IN2(n91), .QN(n55) );
  NOR2X0 U70 ( .IN1(n96), .IN2(n90), .QN(n54) );
  NOR2X0 U71 ( .IN1(n96), .IN2(n89), .QN(n53) );
  NOR2X0 U72 ( .IN1(n92), .IN2(n95), .QN(n51) );
  NOR2X0 U73 ( .IN1(n91), .IN2(n95), .QN(n50) );
  NOR2X0 U74 ( .IN1(n90), .IN2(n95), .QN(n49) );
  NOR2X0 U75 ( .IN1(n89), .IN2(n95), .QN(n48) );
  NOR2X0 U76 ( .IN1(n92), .IN2(n94), .QN(n46) );
  NOR2X0 U77 ( .IN1(n91), .IN2(n94), .QN(n45) );
  NOR2X0 U78 ( .IN1(n90), .IN2(n94), .QN(n44) );
  NOR2X0 U79 ( .IN1(n89), .IN2(n94), .QN(n43) );
  NOR2X0 U80 ( .IN1(n92), .IN2(n93), .QN(n41) );
  NOR2X0 U81 ( .IN1(n91), .IN2(n93), .QN(n40) );
  NOR2X0 U82 ( .IN1(n90), .IN2(n93), .QN(n39) );
  NOR2X0 U83 ( .IN1(n89), .IN2(n93), .QN(n38) );
endmodule


module linear_DW_mult_uns_4 ( a, b, product );
  input [4:0] a;
  input [4:0] b;
  output [9:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n89, n90, n91,
         n92, n93, n94, n95, n96;
  assign n33 = b[3];
  assign n34 = b[2];
  assign n35 = b[1];
  assign n36 = b[0];
  assign n37 = a[3];
  assign n42 = a[2];
  assign n47 = a[1];
  assign n52 = a[0];

  FADDX1 U4 ( .A(n11), .B(n10), .CI(n3), .CO(n2), .S(product[7]) );
  FADDX1 U5 ( .A(n12), .B(n15), .CI(n4), .CO(n3), .S(product[6]) );
  FADDX1 U6 ( .A(n16), .B(n21), .CI(n5), .CO(n4), .S(product[5]) );
  FADDX1 U7 ( .A(n22), .B(n27), .CI(n6), .CO(n5), .S(product[4]) );
  FADDX1 U8 ( .A(n28), .B(n31), .CI(n7), .CO(n6), .S(product[3]) );
  FADDX1 U9 ( .A(n32), .B(n46), .CI(n8), .CO(n7), .S(product[2]) );
  HADDX1 U10 ( .A0(n51), .B0(n55), .C1(n8), .SO(product[1]) );
  FADDX1 U11 ( .A(n33), .B(n37), .CI(n13), .CO(n9), .S(n10) );
  FADDX1 U12 ( .A(n14), .B(n19), .CI(n17), .CO(n11), .S(n12) );
  FADDX1 U13 ( .A(n34), .B(n42), .CI(n38), .CO(n13), .S(n14) );
  FADDX1 U14 ( .A(n23), .B(n25), .CI(n18), .CO(n15), .S(n16) );
  FADDX1 U15 ( .A(n39), .B(n43), .CI(n20), .CO(n17), .S(n18) );
  HADDX1 U16 ( .A0(n47), .B0(n35), .C1(n19), .SO(n20) );
  FADDX1 U17 ( .A(n29), .B(n26), .CI(n24), .CO(n21), .S(n22) );
  FADDX1 U18 ( .A(n40), .B(n48), .CI(n44), .CO(n23), .S(n24) );
  HADDX1 U19 ( .A0(n36), .B0(n52), .C1(n25), .SO(n26) );
  FADDX1 U20 ( .A(n49), .B(n53), .CI(n30), .CO(n27), .S(n28) );
  HADDX1 U21 ( .A0(n45), .B0(n41), .C1(n29), .SO(n30) );
  HADDX1 U22 ( .A0(n54), .B0(n50), .C1(n31), .SO(n32) );
  INVX0 U58 ( .INP(n34), .ZN(n90) );
  INVX0 U59 ( .INP(n42), .ZN(n94) );
  INVX0 U60 ( .INP(n37), .ZN(n93) );
  INVX0 U61 ( .INP(n52), .ZN(n96) );
  INVX0 U62 ( .INP(n47), .ZN(n95) );
  INVX0 U63 ( .INP(n33), .ZN(n89) );
  INVX0 U64 ( .INP(n35), .ZN(n91) );
  INVX0 U65 ( .INP(n36), .ZN(n92) );
  OR2X1 U66 ( .IN1(n2), .IN2(n9), .Q(product[9]) );
  XNOR2X1 U67 ( .IN1(n2), .IN2(n9), .Q(product[8]) );
  NOR2X0 U68 ( .IN1(n96), .IN2(n92), .QN(product[0]) );
  NOR2X0 U69 ( .IN1(n96), .IN2(n91), .QN(n55) );
  NOR2X0 U70 ( .IN1(n96), .IN2(n90), .QN(n54) );
  NOR2X0 U71 ( .IN1(n96), .IN2(n89), .QN(n53) );
  NOR2X0 U72 ( .IN1(n92), .IN2(n95), .QN(n51) );
  NOR2X0 U73 ( .IN1(n91), .IN2(n95), .QN(n50) );
  NOR2X0 U74 ( .IN1(n90), .IN2(n95), .QN(n49) );
  NOR2X0 U75 ( .IN1(n89), .IN2(n95), .QN(n48) );
  NOR2X0 U76 ( .IN1(n92), .IN2(n94), .QN(n46) );
  NOR2X0 U77 ( .IN1(n91), .IN2(n94), .QN(n45) );
  NOR2X0 U78 ( .IN1(n90), .IN2(n94), .QN(n44) );
  NOR2X0 U79 ( .IN1(n89), .IN2(n94), .QN(n43) );
  NOR2X0 U80 ( .IN1(n92), .IN2(n93), .QN(n41) );
  NOR2X0 U81 ( .IN1(n91), .IN2(n93), .QN(n40) );
  NOR2X0 U82 ( .IN1(n90), .IN2(n93), .QN(n39) );
  NOR2X0 U83 ( .IN1(n89), .IN2(n93), .QN(n38) );
endmodule


module linear_DW_mult_uns_5 ( a, b, product );
  input [4:0] a;
  input [4:0] b;
  output [9:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n89, n90, n91,
         n92, n93, n94, n95, n96;
  assign n33 = b[3];
  assign n34 = b[2];
  assign n35 = b[1];
  assign n36 = b[0];
  assign n37 = a[3];
  assign n42 = a[2];
  assign n47 = a[1];
  assign n52 = a[0];

  FADDX1 U4 ( .A(n11), .B(n10), .CI(n3), .CO(n2), .S(product[7]) );
  FADDX1 U5 ( .A(n12), .B(n15), .CI(n4), .CO(n3), .S(product[6]) );
  FADDX1 U6 ( .A(n16), .B(n21), .CI(n5), .CO(n4), .S(product[5]) );
  FADDX1 U7 ( .A(n22), .B(n27), .CI(n6), .CO(n5), .S(product[4]) );
  FADDX1 U8 ( .A(n28), .B(n31), .CI(n7), .CO(n6), .S(product[3]) );
  FADDX1 U9 ( .A(n32), .B(n46), .CI(n8), .CO(n7), .S(product[2]) );
  HADDX1 U10 ( .A0(n51), .B0(n55), .C1(n8), .SO(product[1]) );
  FADDX1 U11 ( .A(n33), .B(n37), .CI(n13), .CO(n9), .S(n10) );
  FADDX1 U12 ( .A(n14), .B(n19), .CI(n17), .CO(n11), .S(n12) );
  FADDX1 U13 ( .A(n34), .B(n42), .CI(n38), .CO(n13), .S(n14) );
  FADDX1 U14 ( .A(n23), .B(n25), .CI(n18), .CO(n15), .S(n16) );
  FADDX1 U15 ( .A(n39), .B(n43), .CI(n20), .CO(n17), .S(n18) );
  HADDX1 U16 ( .A0(n47), .B0(n35), .C1(n19), .SO(n20) );
  FADDX1 U17 ( .A(n29), .B(n26), .CI(n24), .CO(n21), .S(n22) );
  FADDX1 U18 ( .A(n40), .B(n48), .CI(n44), .CO(n23), .S(n24) );
  HADDX1 U19 ( .A0(n36), .B0(n52), .C1(n25), .SO(n26) );
  FADDX1 U20 ( .A(n49), .B(n53), .CI(n30), .CO(n27), .S(n28) );
  HADDX1 U21 ( .A0(n45), .B0(n41), .C1(n29), .SO(n30) );
  HADDX1 U22 ( .A0(n54), .B0(n50), .C1(n31), .SO(n32) );
  INVX0 U58 ( .INP(n34), .ZN(n90) );
  INVX0 U59 ( .INP(n42), .ZN(n94) );
  INVX0 U60 ( .INP(n37), .ZN(n93) );
  INVX0 U61 ( .INP(n52), .ZN(n96) );
  INVX0 U62 ( .INP(n47), .ZN(n95) );
  INVX0 U63 ( .INP(n33), .ZN(n89) );
  INVX0 U64 ( .INP(n35), .ZN(n91) );
  INVX0 U65 ( .INP(n36), .ZN(n92) );
  OR2X1 U66 ( .IN1(n2), .IN2(n9), .Q(product[9]) );
  XNOR2X1 U67 ( .IN1(n2), .IN2(n9), .Q(product[8]) );
  NOR2X0 U68 ( .IN1(n96), .IN2(n92), .QN(product[0]) );
  NOR2X0 U69 ( .IN1(n96), .IN2(n91), .QN(n55) );
  NOR2X0 U70 ( .IN1(n96), .IN2(n90), .QN(n54) );
  NOR2X0 U71 ( .IN1(n96), .IN2(n89), .QN(n53) );
  NOR2X0 U72 ( .IN1(n92), .IN2(n95), .QN(n51) );
  NOR2X0 U73 ( .IN1(n91), .IN2(n95), .QN(n50) );
  NOR2X0 U74 ( .IN1(n90), .IN2(n95), .QN(n49) );
  NOR2X0 U75 ( .IN1(n89), .IN2(n95), .QN(n48) );
  NOR2X0 U76 ( .IN1(n92), .IN2(n94), .QN(n46) );
  NOR2X0 U77 ( .IN1(n91), .IN2(n94), .QN(n45) );
  NOR2X0 U78 ( .IN1(n90), .IN2(n94), .QN(n44) );
  NOR2X0 U79 ( .IN1(n89), .IN2(n94), .QN(n43) );
  NOR2X0 U80 ( .IN1(n92), .IN2(n93), .QN(n41) );
  NOR2X0 U81 ( .IN1(n91), .IN2(n93), .QN(n40) );
  NOR2X0 U82 ( .IN1(n90), .IN2(n93), .QN(n39) );
  NOR2X0 U83 ( .IN1(n89), .IN2(n93), .QN(n38) );
endmodule


module linear_DW_mult_uns_6 ( a, b, product );
  input [4:0] a;
  input [4:0] b;
  output [9:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n89, n90, n91,
         n92, n93, n94, n95, n96;
  assign n33 = b[3];
  assign n34 = b[2];
  assign n35 = b[1];
  assign n36 = b[0];
  assign n37 = a[3];
  assign n42 = a[2];
  assign n47 = a[1];
  assign n52 = a[0];

  FADDX1 U4 ( .A(n11), .B(n10), .CI(n3), .CO(n2), .S(product[7]) );
  FADDX1 U5 ( .A(n12), .B(n15), .CI(n4), .CO(n3), .S(product[6]) );
  FADDX1 U6 ( .A(n16), .B(n21), .CI(n5), .CO(n4), .S(product[5]) );
  FADDX1 U7 ( .A(n22), .B(n27), .CI(n6), .CO(n5), .S(product[4]) );
  FADDX1 U8 ( .A(n28), .B(n31), .CI(n7), .CO(n6), .S(product[3]) );
  FADDX1 U9 ( .A(n32), .B(n46), .CI(n8), .CO(n7), .S(product[2]) );
  HADDX1 U10 ( .A0(n51), .B0(n55), .C1(n8), .SO(product[1]) );
  FADDX1 U11 ( .A(n33), .B(n37), .CI(n13), .CO(n9), .S(n10) );
  FADDX1 U12 ( .A(n14), .B(n19), .CI(n17), .CO(n11), .S(n12) );
  FADDX1 U13 ( .A(n34), .B(n42), .CI(n38), .CO(n13), .S(n14) );
  FADDX1 U14 ( .A(n23), .B(n25), .CI(n18), .CO(n15), .S(n16) );
  FADDX1 U15 ( .A(n39), .B(n43), .CI(n20), .CO(n17), .S(n18) );
  HADDX1 U16 ( .A0(n47), .B0(n35), .C1(n19), .SO(n20) );
  FADDX1 U17 ( .A(n29), .B(n26), .CI(n24), .CO(n21), .S(n22) );
  FADDX1 U18 ( .A(n40), .B(n48), .CI(n44), .CO(n23), .S(n24) );
  HADDX1 U19 ( .A0(n36), .B0(n52), .C1(n25), .SO(n26) );
  FADDX1 U20 ( .A(n49), .B(n53), .CI(n30), .CO(n27), .S(n28) );
  HADDX1 U21 ( .A0(n45), .B0(n41), .C1(n29), .SO(n30) );
  HADDX1 U22 ( .A0(n54), .B0(n50), .C1(n31), .SO(n32) );
  INVX0 U58 ( .INP(n34), .ZN(n90) );
  INVX0 U59 ( .INP(n42), .ZN(n94) );
  INVX0 U60 ( .INP(n37), .ZN(n93) );
  INVX0 U61 ( .INP(n52), .ZN(n96) );
  INVX0 U62 ( .INP(n47), .ZN(n95) );
  INVX0 U63 ( .INP(n33), .ZN(n89) );
  INVX0 U64 ( .INP(n35), .ZN(n91) );
  INVX0 U65 ( .INP(n36), .ZN(n92) );
  OR2X1 U66 ( .IN1(n2), .IN2(n9), .Q(product[9]) );
  XNOR2X1 U67 ( .IN1(n2), .IN2(n9), .Q(product[8]) );
  NOR2X0 U68 ( .IN1(n96), .IN2(n92), .QN(product[0]) );
  NOR2X0 U69 ( .IN1(n96), .IN2(n91), .QN(n55) );
  NOR2X0 U70 ( .IN1(n96), .IN2(n90), .QN(n54) );
  NOR2X0 U71 ( .IN1(n96), .IN2(n89), .QN(n53) );
  NOR2X0 U72 ( .IN1(n92), .IN2(n95), .QN(n51) );
  NOR2X0 U73 ( .IN1(n91), .IN2(n95), .QN(n50) );
  NOR2X0 U74 ( .IN1(n90), .IN2(n95), .QN(n49) );
  NOR2X0 U75 ( .IN1(n89), .IN2(n95), .QN(n48) );
  NOR2X0 U76 ( .IN1(n92), .IN2(n94), .QN(n46) );
  NOR2X0 U77 ( .IN1(n91), .IN2(n94), .QN(n45) );
  NOR2X0 U78 ( .IN1(n90), .IN2(n94), .QN(n44) );
  NOR2X0 U79 ( .IN1(n89), .IN2(n94), .QN(n43) );
  NOR2X0 U80 ( .IN1(n92), .IN2(n93), .QN(n41) );
  NOR2X0 U81 ( .IN1(n91), .IN2(n93), .QN(n40) );
  NOR2X0 U82 ( .IN1(n90), .IN2(n93), .QN(n39) );
  NOR2X0 U83 ( .IN1(n89), .IN2(n93), .QN(n38) );
endmodule


module linear_DW_mult_uns_7 ( a, b, product );
  input [4:0] a;
  input [4:0] b;
  output [9:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n89, n90, n91,
         n92, n93, n94, n95, n96;
  assign n33 = b[3];
  assign n34 = b[2];
  assign n35 = b[1];
  assign n36 = b[0];
  assign n37 = a[3];
  assign n42 = a[2];
  assign n47 = a[1];
  assign n52 = a[0];

  FADDX1 U4 ( .A(n11), .B(n10), .CI(n3), .CO(n2), .S(product[7]) );
  FADDX1 U5 ( .A(n12), .B(n15), .CI(n4), .CO(n3), .S(product[6]) );
  FADDX1 U6 ( .A(n16), .B(n21), .CI(n5), .CO(n4), .S(product[5]) );
  FADDX1 U7 ( .A(n22), .B(n27), .CI(n6), .CO(n5), .S(product[4]) );
  FADDX1 U8 ( .A(n28), .B(n31), .CI(n7), .CO(n6), .S(product[3]) );
  FADDX1 U9 ( .A(n32), .B(n46), .CI(n8), .CO(n7), .S(product[2]) );
  HADDX1 U10 ( .A0(n51), .B0(n55), .C1(n8), .SO(product[1]) );
  FADDX1 U11 ( .A(n33), .B(n37), .CI(n13), .CO(n9), .S(n10) );
  FADDX1 U12 ( .A(n14), .B(n19), .CI(n17), .CO(n11), .S(n12) );
  FADDX1 U13 ( .A(n34), .B(n42), .CI(n38), .CO(n13), .S(n14) );
  FADDX1 U14 ( .A(n23), .B(n25), .CI(n18), .CO(n15), .S(n16) );
  FADDX1 U15 ( .A(n39), .B(n43), .CI(n20), .CO(n17), .S(n18) );
  HADDX1 U16 ( .A0(n47), .B0(n35), .C1(n19), .SO(n20) );
  FADDX1 U17 ( .A(n29), .B(n26), .CI(n24), .CO(n21), .S(n22) );
  FADDX1 U18 ( .A(n40), .B(n48), .CI(n44), .CO(n23), .S(n24) );
  HADDX1 U19 ( .A0(n36), .B0(n52), .C1(n25), .SO(n26) );
  FADDX1 U20 ( .A(n49), .B(n53), .CI(n30), .CO(n27), .S(n28) );
  HADDX1 U21 ( .A0(n45), .B0(n41), .C1(n29), .SO(n30) );
  HADDX1 U22 ( .A0(n54), .B0(n50), .C1(n31), .SO(n32) );
  INVX0 U58 ( .INP(n34), .ZN(n90) );
  INVX0 U59 ( .INP(n42), .ZN(n94) );
  INVX0 U60 ( .INP(n37), .ZN(n93) );
  INVX0 U61 ( .INP(n52), .ZN(n96) );
  INVX0 U62 ( .INP(n47), .ZN(n95) );
  INVX0 U63 ( .INP(n33), .ZN(n89) );
  INVX0 U64 ( .INP(n35), .ZN(n91) );
  INVX0 U65 ( .INP(n36), .ZN(n92) );
  OR2X1 U66 ( .IN1(n2), .IN2(n9), .Q(product[9]) );
  XNOR2X1 U67 ( .IN1(n2), .IN2(n9), .Q(product[8]) );
  NOR2X0 U68 ( .IN1(n96), .IN2(n92), .QN(product[0]) );
  NOR2X0 U69 ( .IN1(n96), .IN2(n91), .QN(n55) );
  NOR2X0 U70 ( .IN1(n96), .IN2(n90), .QN(n54) );
  NOR2X0 U71 ( .IN1(n96), .IN2(n89), .QN(n53) );
  NOR2X0 U72 ( .IN1(n92), .IN2(n95), .QN(n51) );
  NOR2X0 U73 ( .IN1(n91), .IN2(n95), .QN(n50) );
  NOR2X0 U74 ( .IN1(n90), .IN2(n95), .QN(n49) );
  NOR2X0 U75 ( .IN1(n89), .IN2(n95), .QN(n48) );
  NOR2X0 U76 ( .IN1(n92), .IN2(n94), .QN(n46) );
  NOR2X0 U77 ( .IN1(n91), .IN2(n94), .QN(n45) );
  NOR2X0 U78 ( .IN1(n90), .IN2(n94), .QN(n44) );
  NOR2X0 U79 ( .IN1(n89), .IN2(n94), .QN(n43) );
  NOR2X0 U80 ( .IN1(n92), .IN2(n93), .QN(n41) );
  NOR2X0 U81 ( .IN1(n91), .IN2(n93), .QN(n40) );
  NOR2X0 U82 ( .IN1(n90), .IN2(n93), .QN(n39) );
  NOR2X0 U83 ( .IN1(n89), .IN2(n93), .QN(n38) );
endmodule


module linear_DW_mult_uns_8 ( a, b, product );
  input [4:0] a;
  input [4:0] b;
  output [9:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n89, n90, n91,
         n92, n93, n94, n95, n96;
  assign n33 = b[3];
  assign n34 = b[2];
  assign n35 = b[1];
  assign n36 = b[0];
  assign n37 = a[3];
  assign n42 = a[2];
  assign n47 = a[1];
  assign n52 = a[0];

  FADDX1 U4 ( .A(n11), .B(n10), .CI(n3), .CO(n2), .S(product[7]) );
  FADDX1 U5 ( .A(n12), .B(n15), .CI(n4), .CO(n3), .S(product[6]) );
  FADDX1 U6 ( .A(n16), .B(n21), .CI(n5), .CO(n4), .S(product[5]) );
  FADDX1 U7 ( .A(n22), .B(n27), .CI(n6), .CO(n5), .S(product[4]) );
  FADDX1 U8 ( .A(n28), .B(n31), .CI(n7), .CO(n6), .S(product[3]) );
  FADDX1 U9 ( .A(n32), .B(n46), .CI(n8), .CO(n7), .S(product[2]) );
  HADDX1 U10 ( .A0(n51), .B0(n55), .C1(n8), .SO(product[1]) );
  FADDX1 U11 ( .A(n33), .B(n37), .CI(n13), .CO(n9), .S(n10) );
  FADDX1 U12 ( .A(n14), .B(n19), .CI(n17), .CO(n11), .S(n12) );
  FADDX1 U13 ( .A(n34), .B(n42), .CI(n38), .CO(n13), .S(n14) );
  FADDX1 U14 ( .A(n23), .B(n25), .CI(n18), .CO(n15), .S(n16) );
  FADDX1 U15 ( .A(n39), .B(n43), .CI(n20), .CO(n17), .S(n18) );
  HADDX1 U16 ( .A0(n47), .B0(n35), .C1(n19), .SO(n20) );
  FADDX1 U17 ( .A(n29), .B(n26), .CI(n24), .CO(n21), .S(n22) );
  FADDX1 U18 ( .A(n40), .B(n48), .CI(n44), .CO(n23), .S(n24) );
  HADDX1 U19 ( .A0(n36), .B0(n52), .C1(n25), .SO(n26) );
  FADDX1 U20 ( .A(n49), .B(n53), .CI(n30), .CO(n27), .S(n28) );
  HADDX1 U21 ( .A0(n45), .B0(n41), .C1(n29), .SO(n30) );
  HADDX1 U22 ( .A0(n54), .B0(n50), .C1(n31), .SO(n32) );
  INVX0 U58 ( .INP(n34), .ZN(n90) );
  INVX0 U59 ( .INP(n42), .ZN(n94) );
  INVX0 U60 ( .INP(n37), .ZN(n93) );
  INVX0 U61 ( .INP(n52), .ZN(n96) );
  INVX0 U62 ( .INP(n47), .ZN(n95) );
  INVX0 U63 ( .INP(n33), .ZN(n89) );
  INVX0 U64 ( .INP(n35), .ZN(n91) );
  INVX0 U65 ( .INP(n36), .ZN(n92) );
  OR2X1 U66 ( .IN1(n2), .IN2(n9), .Q(product[9]) );
  XNOR2X1 U67 ( .IN1(n2), .IN2(n9), .Q(product[8]) );
  NOR2X0 U68 ( .IN1(n96), .IN2(n92), .QN(product[0]) );
  NOR2X0 U69 ( .IN1(n96), .IN2(n91), .QN(n55) );
  NOR2X0 U70 ( .IN1(n96), .IN2(n90), .QN(n54) );
  NOR2X0 U71 ( .IN1(n96), .IN2(n89), .QN(n53) );
  NOR2X0 U72 ( .IN1(n92), .IN2(n95), .QN(n51) );
  NOR2X0 U73 ( .IN1(n91), .IN2(n95), .QN(n50) );
  NOR2X0 U74 ( .IN1(n90), .IN2(n95), .QN(n49) );
  NOR2X0 U75 ( .IN1(n89), .IN2(n95), .QN(n48) );
  NOR2X0 U76 ( .IN1(n92), .IN2(n94), .QN(n46) );
  NOR2X0 U77 ( .IN1(n91), .IN2(n94), .QN(n45) );
  NOR2X0 U78 ( .IN1(n90), .IN2(n94), .QN(n44) );
  NOR2X0 U79 ( .IN1(n89), .IN2(n94), .QN(n43) );
  NOR2X0 U80 ( .IN1(n92), .IN2(n93), .QN(n41) );
  NOR2X0 U81 ( .IN1(n91), .IN2(n93), .QN(n40) );
  NOR2X0 U82 ( .IN1(n90), .IN2(n93), .QN(n39) );
  NOR2X0 U83 ( .IN1(n89), .IN2(n93), .QN(n38) );
endmodule


module linear_DW_mult_uns_9 ( a, b, product );
  input [4:0] a;
  input [4:0] b;
  output [9:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n89, n90, n91,
         n92, n93, n94, n95, n96;
  assign n33 = b[3];
  assign n34 = b[2];
  assign n35 = b[1];
  assign n36 = b[0];
  assign n37 = a[3];
  assign n42 = a[2];
  assign n47 = a[1];
  assign n52 = a[0];

  FADDX1 U4 ( .A(n11), .B(n10), .CI(n3), .CO(n2), .S(product[7]) );
  FADDX1 U5 ( .A(n12), .B(n15), .CI(n4), .CO(n3), .S(product[6]) );
  FADDX1 U6 ( .A(n16), .B(n21), .CI(n5), .CO(n4), .S(product[5]) );
  FADDX1 U7 ( .A(n22), .B(n27), .CI(n6), .CO(n5), .S(product[4]) );
  FADDX1 U8 ( .A(n28), .B(n31), .CI(n7), .CO(n6), .S(product[3]) );
  FADDX1 U9 ( .A(n32), .B(n46), .CI(n8), .CO(n7), .S(product[2]) );
  HADDX1 U10 ( .A0(n51), .B0(n55), .C1(n8), .SO(product[1]) );
  FADDX1 U11 ( .A(n33), .B(n37), .CI(n13), .CO(n9), .S(n10) );
  FADDX1 U12 ( .A(n14), .B(n19), .CI(n17), .CO(n11), .S(n12) );
  FADDX1 U13 ( .A(n34), .B(n42), .CI(n38), .CO(n13), .S(n14) );
  FADDX1 U14 ( .A(n23), .B(n25), .CI(n18), .CO(n15), .S(n16) );
  FADDX1 U15 ( .A(n39), .B(n43), .CI(n20), .CO(n17), .S(n18) );
  HADDX1 U16 ( .A0(n47), .B0(n35), .C1(n19), .SO(n20) );
  FADDX1 U17 ( .A(n29), .B(n26), .CI(n24), .CO(n21), .S(n22) );
  FADDX1 U18 ( .A(n40), .B(n48), .CI(n44), .CO(n23), .S(n24) );
  HADDX1 U19 ( .A0(n36), .B0(n52), .C1(n25), .SO(n26) );
  FADDX1 U20 ( .A(n49), .B(n53), .CI(n30), .CO(n27), .S(n28) );
  HADDX1 U21 ( .A0(n45), .B0(n41), .C1(n29), .SO(n30) );
  HADDX1 U22 ( .A0(n54), .B0(n50), .C1(n31), .SO(n32) );
  INVX0 U58 ( .INP(n34), .ZN(n90) );
  INVX0 U59 ( .INP(n42), .ZN(n94) );
  INVX0 U60 ( .INP(n37), .ZN(n93) );
  INVX0 U61 ( .INP(n52), .ZN(n96) );
  INVX0 U62 ( .INP(n47), .ZN(n95) );
  INVX0 U63 ( .INP(n33), .ZN(n89) );
  INVX0 U64 ( .INP(n35), .ZN(n91) );
  INVX0 U65 ( .INP(n36), .ZN(n92) );
  OR2X1 U66 ( .IN1(n2), .IN2(n9), .Q(product[9]) );
  XNOR2X1 U67 ( .IN1(n2), .IN2(n9), .Q(product[8]) );
  NOR2X0 U68 ( .IN1(n96), .IN2(n92), .QN(product[0]) );
  NOR2X0 U69 ( .IN1(n96), .IN2(n91), .QN(n55) );
  NOR2X0 U70 ( .IN1(n96), .IN2(n90), .QN(n54) );
  NOR2X0 U71 ( .IN1(n96), .IN2(n89), .QN(n53) );
  NOR2X0 U72 ( .IN1(n92), .IN2(n95), .QN(n51) );
  NOR2X0 U73 ( .IN1(n91), .IN2(n95), .QN(n50) );
  NOR2X0 U74 ( .IN1(n90), .IN2(n95), .QN(n49) );
  NOR2X0 U75 ( .IN1(n89), .IN2(n95), .QN(n48) );
  NOR2X0 U76 ( .IN1(n92), .IN2(n94), .QN(n46) );
  NOR2X0 U77 ( .IN1(n91), .IN2(n94), .QN(n45) );
  NOR2X0 U78 ( .IN1(n90), .IN2(n94), .QN(n44) );
  NOR2X0 U79 ( .IN1(n89), .IN2(n94), .QN(n43) );
  NOR2X0 U80 ( .IN1(n92), .IN2(n93), .QN(n41) );
  NOR2X0 U81 ( .IN1(n91), .IN2(n93), .QN(n40) );
  NOR2X0 U82 ( .IN1(n90), .IN2(n93), .QN(n39) );
  NOR2X0 U83 ( .IN1(n89), .IN2(n93), .QN(n38) );
endmodule


module linear ( clk, rst, p__arg0_0_0, p__arg0_0_1, p__arg0_0_10, p__arg0_0_2, 
        p__arg0_0_3, p__arg0_0_4, p__arg0_0_5, p__arg0_0_6, p__arg0_0_7, 
        p__arg0_0_8, p__arg0_0_9, p___constant_11x11xf32_0_0, 
        p___constant_11x11xf32_0_1, p___constant_11x11xf32_0_10, 
        p___constant_11x11xf32_0_2, p___constant_11x11xf32_0_3, 
        p___constant_11x11xf32_0_4, p___constant_11x11xf32_0_5, 
        p___constant_11x11xf32_0_6, p___constant_11x11xf32_0_7, 
        p___constant_11x11xf32_0_8, p___constant_11x11xf32_0_9, 
        p___constant_11x11xf32_10_0, p___constant_11x11xf32_10_1, 
        p___constant_11x11xf32_10_10, p___constant_11x11xf32_10_2, 
        p___constant_11x11xf32_10_3, p___constant_11x11xf32_10_4, 
        p___constant_11x11xf32_10_5, p___constant_11x11xf32_10_6, 
        p___constant_11x11xf32_10_7, p___constant_11x11xf32_10_8, 
        p___constant_11x11xf32_10_9, p___constant_11x11xf32_1_0, 
        p___constant_11x11xf32_1_1, p___constant_11x11xf32_1_10, 
        p___constant_11x11xf32_1_2, p___constant_11x11xf32_1_3, 
        p___constant_11x11xf32_1_4, p___constant_11x11xf32_1_5, 
        p___constant_11x11xf32_1_6, p___constant_11x11xf32_1_7, 
        p___constant_11x11xf32_1_8, p___constant_11x11xf32_1_9, 
        p___constant_11x11xf32_2_0, p___constant_11x11xf32_2_1, 
        p___constant_11x11xf32_2_10, p___constant_11x11xf32_2_2, 
        p___constant_11x11xf32_2_3, p___constant_11x11xf32_2_4, 
        p___constant_11x11xf32_2_5, p___constant_11x11xf32_2_6, 
        p___constant_11x11xf32_2_7, p___constant_11x11xf32_2_8, 
        p___constant_11x11xf32_2_9, p___constant_11x11xf32_3_0, 
        p___constant_11x11xf32_3_1, p___constant_11x11xf32_3_10, 
        p___constant_11x11xf32_3_2, p___constant_11x11xf32_3_3, 
        p___constant_11x11xf32_3_4, p___constant_11x11xf32_3_5, 
        p___constant_11x11xf32_3_6, p___constant_11x11xf32_3_7, 
        p___constant_11x11xf32_3_8, p___constant_11x11xf32_3_9, 
        p___constant_11x11xf32_4_0, p___constant_11x11xf32_4_1, 
        p___constant_11x11xf32_4_10, p___constant_11x11xf32_4_2, 
        p___constant_11x11xf32_4_3, p___constant_11x11xf32_4_4, 
        p___constant_11x11xf32_4_5, p___constant_11x11xf32_4_6, 
        p___constant_11x11xf32_4_7, p___constant_11x11xf32_4_8, 
        p___constant_11x11xf32_4_9, p___constant_11x11xf32_5_0, 
        p___constant_11x11xf32_5_1, p___constant_11x11xf32_5_10, 
        p___constant_11x11xf32_5_2, p___constant_11x11xf32_5_3, 
        p___constant_11x11xf32_5_4, p___constant_11x11xf32_5_5, 
        p___constant_11x11xf32_5_6, p___constant_11x11xf32_5_7, 
        p___constant_11x11xf32_5_8, p___constant_11x11xf32_5_9, 
        p___constant_11x11xf32_6_0, p___constant_11x11xf32_6_1, 
        p___constant_11x11xf32_6_10, p___constant_11x11xf32_6_2, 
        p___constant_11x11xf32_6_3, p___constant_11x11xf32_6_4, 
        p___constant_11x11xf32_6_5, p___constant_11x11xf32_6_6, 
        p___constant_11x11xf32_6_7, p___constant_11x11xf32_6_8, 
        p___constant_11x11xf32_6_9, p___constant_11x11xf32_7_0, 
        p___constant_11x11xf32_7_1, p___constant_11x11xf32_7_10, 
        p___constant_11x11xf32_7_2, p___constant_11x11xf32_7_3, 
        p___constant_11x11xf32_7_4, p___constant_11x11xf32_7_5, 
        p___constant_11x11xf32_7_6, p___constant_11x11xf32_7_7, 
        p___constant_11x11xf32_7_8, p___constant_11x11xf32_7_9, 
        p___constant_11x11xf32_8_0, p___constant_11x11xf32_8_1, 
        p___constant_11x11xf32_8_10, p___constant_11x11xf32_8_2, 
        p___constant_11x11xf32_8_3, p___constant_11x11xf32_8_4, 
        p___constant_11x11xf32_8_5, p___constant_11x11xf32_8_6, 
        p___constant_11x11xf32_8_7, p___constant_11x11xf32_8_8, 
        p___constant_11x11xf32_8_9, p___constant_11x11xf32_9_0, 
        p___constant_11x11xf32_9_1, p___constant_11x11xf32_9_10, 
        p___constant_11x11xf32_9_2, p___constant_11x11xf32_9_3, 
        p___constant_11x11xf32_9_4, p___constant_11x11xf32_9_5, 
        p___constant_11x11xf32_9_6, p___constant_11x11xf32_9_7, 
        p___constant_11x11xf32_9_8, p___constant_11x11xf32_9_9, 
        p___constant_11xf32_0, p___constant_11xf32_1, p___constant_11xf32_10, 
        p___constant_11xf32_2, p___constant_11xf32_3, p___constant_11xf32_4, 
        p___constant_11xf32_5, p___constant_11xf32_6, p___constant_11xf32_7, 
        p___constant_11xf32_8, p___constant_11xf32_9, output_p_val_313 );
  input [11:0] p__arg0_0_0;
  input [11:0] p__arg0_0_1;
  input [11:0] p__arg0_0_10;
  input [11:0] p__arg0_0_2;
  input [11:0] p__arg0_0_3;
  input [11:0] p__arg0_0_4;
  input [11:0] p__arg0_0_5;
  input [11:0] p__arg0_0_6;
  input [11:0] p__arg0_0_7;
  input [11:0] p__arg0_0_8;
  input [11:0] p__arg0_0_9;
  input [11:0] p___constant_11x11xf32_0_0;
  input [11:0] p___constant_11x11xf32_0_1;
  input [11:0] p___constant_11x11xf32_0_10;
  input [11:0] p___constant_11x11xf32_0_2;
  input [11:0] p___constant_11x11xf32_0_3;
  input [11:0] p___constant_11x11xf32_0_4;
  input [11:0] p___constant_11x11xf32_0_5;
  input [11:0] p___constant_11x11xf32_0_6;
  input [11:0] p___constant_11x11xf32_0_7;
  input [11:0] p___constant_11x11xf32_0_8;
  input [11:0] p___constant_11x11xf32_0_9;
  input [11:0] p___constant_11x11xf32_10_0;
  input [11:0] p___constant_11x11xf32_10_1;
  input [11:0] p___constant_11x11xf32_10_10;
  input [11:0] p___constant_11x11xf32_10_2;
  input [11:0] p___constant_11x11xf32_10_3;
  input [11:0] p___constant_11x11xf32_10_4;
  input [11:0] p___constant_11x11xf32_10_5;
  input [11:0] p___constant_11x11xf32_10_6;
  input [11:0] p___constant_11x11xf32_10_7;
  input [11:0] p___constant_11x11xf32_10_8;
  input [11:0] p___constant_11x11xf32_10_9;
  input [11:0] p___constant_11x11xf32_1_0;
  input [11:0] p___constant_11x11xf32_1_1;
  input [11:0] p___constant_11x11xf32_1_10;
  input [11:0] p___constant_11x11xf32_1_2;
  input [11:0] p___constant_11x11xf32_1_3;
  input [11:0] p___constant_11x11xf32_1_4;
  input [11:0] p___constant_11x11xf32_1_5;
  input [11:0] p___constant_11x11xf32_1_6;
  input [11:0] p___constant_11x11xf32_1_7;
  input [11:0] p___constant_11x11xf32_1_8;
  input [11:0] p___constant_11x11xf32_1_9;
  input [11:0] p___constant_11x11xf32_2_0;
  input [11:0] p___constant_11x11xf32_2_1;
  input [11:0] p___constant_11x11xf32_2_10;
  input [11:0] p___constant_11x11xf32_2_2;
  input [11:0] p___constant_11x11xf32_2_3;
  input [11:0] p___constant_11x11xf32_2_4;
  input [11:0] p___constant_11x11xf32_2_5;
  input [11:0] p___constant_11x11xf32_2_6;
  input [11:0] p___constant_11x11xf32_2_7;
  input [11:0] p___constant_11x11xf32_2_8;
  input [11:0] p___constant_11x11xf32_2_9;
  input [11:0] p___constant_11x11xf32_3_0;
  input [11:0] p___constant_11x11xf32_3_1;
  input [11:0] p___constant_11x11xf32_3_10;
  input [11:0] p___constant_11x11xf32_3_2;
  input [11:0] p___constant_11x11xf32_3_3;
  input [11:0] p___constant_11x11xf32_3_4;
  input [11:0] p___constant_11x11xf32_3_5;
  input [11:0] p___constant_11x11xf32_3_6;
  input [11:0] p___constant_11x11xf32_3_7;
  input [11:0] p___constant_11x11xf32_3_8;
  input [11:0] p___constant_11x11xf32_3_9;
  input [11:0] p___constant_11x11xf32_4_0;
  input [11:0] p___constant_11x11xf32_4_1;
  input [11:0] p___constant_11x11xf32_4_10;
  input [11:0] p___constant_11x11xf32_4_2;
  input [11:0] p___constant_11x11xf32_4_3;
  input [11:0] p___constant_11x11xf32_4_4;
  input [11:0] p___constant_11x11xf32_4_5;
  input [11:0] p___constant_11x11xf32_4_6;
  input [11:0] p___constant_11x11xf32_4_7;
  input [11:0] p___constant_11x11xf32_4_8;
  input [11:0] p___constant_11x11xf32_4_9;
  input [11:0] p___constant_11x11xf32_5_0;
  input [11:0] p___constant_11x11xf32_5_1;
  input [11:0] p___constant_11x11xf32_5_10;
  input [11:0] p___constant_11x11xf32_5_2;
  input [11:0] p___constant_11x11xf32_5_3;
  input [11:0] p___constant_11x11xf32_5_4;
  input [11:0] p___constant_11x11xf32_5_5;
  input [11:0] p___constant_11x11xf32_5_6;
  input [11:0] p___constant_11x11xf32_5_7;
  input [11:0] p___constant_11x11xf32_5_8;
  input [11:0] p___constant_11x11xf32_5_9;
  input [11:0] p___constant_11x11xf32_6_0;
  input [11:0] p___constant_11x11xf32_6_1;
  input [11:0] p___constant_11x11xf32_6_10;
  input [11:0] p___constant_11x11xf32_6_2;
  input [11:0] p___constant_11x11xf32_6_3;
  input [11:0] p___constant_11x11xf32_6_4;
  input [11:0] p___constant_11x11xf32_6_5;
  input [11:0] p___constant_11x11xf32_6_6;
  input [11:0] p___constant_11x11xf32_6_7;
  input [11:0] p___constant_11x11xf32_6_8;
  input [11:0] p___constant_11x11xf32_6_9;
  input [11:0] p___constant_11x11xf32_7_0;
  input [11:0] p___constant_11x11xf32_7_1;
  input [11:0] p___constant_11x11xf32_7_10;
  input [11:0] p___constant_11x11xf32_7_2;
  input [11:0] p___constant_11x11xf32_7_3;
  input [11:0] p___constant_11x11xf32_7_4;
  input [11:0] p___constant_11x11xf32_7_5;
  input [11:0] p___constant_11x11xf32_7_6;
  input [11:0] p___constant_11x11xf32_7_7;
  input [11:0] p___constant_11x11xf32_7_8;
  input [11:0] p___constant_11x11xf32_7_9;
  input [11:0] p___constant_11x11xf32_8_0;
  input [11:0] p___constant_11x11xf32_8_1;
  input [11:0] p___constant_11x11xf32_8_10;
  input [11:0] p___constant_11x11xf32_8_2;
  input [11:0] p___constant_11x11xf32_8_3;
  input [11:0] p___constant_11x11xf32_8_4;
  input [11:0] p___constant_11x11xf32_8_5;
  input [11:0] p___constant_11x11xf32_8_6;
  input [11:0] p___constant_11x11xf32_8_7;
  input [11:0] p___constant_11x11xf32_8_8;
  input [11:0] p___constant_11x11xf32_8_9;
  input [11:0] p___constant_11x11xf32_9_0;
  input [11:0] p___constant_11x11xf32_9_1;
  input [11:0] p___constant_11x11xf32_9_10;
  input [11:0] p___constant_11x11xf32_9_2;
  input [11:0] p___constant_11x11xf32_9_3;
  input [11:0] p___constant_11x11xf32_9_4;
  input [11:0] p___constant_11x11xf32_9_5;
  input [11:0] p___constant_11x11xf32_9_6;
  input [11:0] p___constant_11x11xf32_9_7;
  input [11:0] p___constant_11x11xf32_9_8;
  input [11:0] p___constant_11x11xf32_9_9;
  input [11:0] p___constant_11xf32_0;
  input [11:0] p___constant_11xf32_1;
  input [11:0] p___constant_11xf32_10;
  input [11:0] p___constant_11xf32_2;
  input [11:0] p___constant_11xf32_3;
  input [11:0] p___constant_11xf32_4;
  input [11:0] p___constant_11xf32_5;
  input [11:0] p___constant_11xf32_6;
  input [11:0] p___constant_11xf32_7;
  input [11:0] p___constant_11xf32_8;
  input [11:0] p___constant_11xf32_9;
  output [11:0] output_p_val_313;
  input clk, rst;
  wire   n5302, n5301, n5300, n5299, n5298, n5297, n5296, n5295, n5294, n5314,
         n5313, n5312, n5311, n5310, n5309, n5308, n5307, n5306, n5338, n5337,
         n5336, n5335, n5334, n5350, n5349, n5348, n5347, n5346, n5374, n5373,
         n5372, n5371, n5370, n5369, n5368, n5367, n5366, n5386, n5385, n5384,
         n5383, n5382, n5381, n5380, n5379, n5378, n5410, n5409, n5408, n5407,
         n5406, n5422, n5421, n5420, n5419, n5418, n5446, n5445, n5444, n5443,
         n5442, n5441, n5440, n5439, n5438, n5458, n5457, n5456, n5455, n5454,
         n5453, n5452, n5451, n5450, n5482, n5481, n5480, n5479, n5478, n5494,
         n5493, n5492, n5491, n5490, n5518, n5517, n5516, n5515, n5514, n5513,
         n5512, n5511, n5510, n5530, n5529, n5528, n5527, n5526, n5525, n5524,
         n5523, n5522, n5554, n5553, n5552, n5551, n5550, n5566, n5565, n5564,
         n5563, n5562, n5590, n5589, n5588, n5587, n5586, n5585, n5584, n5583,
         n5582, n5602, n5601, n5600, n5599, n5598, n5597, n5596, n5595, n5594,
         n5626, n5625, n5624, n5623, n5622, n5638, n5637, n5636, n5635, n5634,
         n5662, n5661, n5660, n5659, n5658, n5657, n5656, n5655, n5654, n5674,
         n5673, n5672, n5671, n5670, n5669, n5668, n5667, n5666, n5698, n5697,
         n5696, n5695, n5694, n5710, n5709, n5708, n5707, n5706, n5734, n5733,
         n5732, n5731, n5730, n5729, n5728, n5727, n5726, n5746, n5745, n5744,
         n5743, n5742, n5741, n5740, n5739, n5738, n5770, n5769, n5768, n5767,
         n5766, n5782, n5781, n5780, n5779, n5778, n5806, n5805, n5804, n5803,
         n5802, n5801, n5800, n5799, n5798, n5818, n5817, n5816, n5815, n5814,
         n5813, n5812, n5811, n5810, n5842, n5841, n5840, n5839, n5838, n5854,
         n5853, n5852, n5851, n5850, n5878, n5877, n5876, n5875, n5874, n5873,
         n5872, n5871, n5870, n5890, n5889, n5888, n5887, n5886, n5885, n5884,
         n5883, n5882, n5914, n5913, n5912, n5911, n5910, n5926, n5925, n5924,
         n5923, n5922, n5950, n5949, n5948, n5947, n5946, n5945, n5944, n5943,
         n5942, n5962, n5961, n5960, n5959, n5958, n5957, n5956, n5955, n5954,
         n5986, n5985, n5984, n5983, n5982, n5998, n5997, n5996, n5995, n5994,
         \U616/DATA2_0 , \U616/DATA2_1 , \U616/DATA2_2 , \U616/DATA2_3 ,
         \U616/DATA2_4 , \U616/DATA2_5 , \U616/DATA2_6 , \U616/DATA2_7 ,
         \U616/DATA2_8 , \U616/DATA2_9 , \U616/DATA2_10 , \U616/DATA2_11 ,
         \U616/DATA1_0 , \U616/DATA1_1 , \U616/DATA1_2 , \U616/DATA1_3 ,
         \U616/DATA1_4 , \U616/DATA1_5 , \U616/DATA1_6 , \U616/DATA1_7 ,
         \U616/DATA1_8 , \U616/DATA1_9 , \U616/DATA1_10 , \U616/DATA1_11 ,
         \U615/DATA2_0 , \U615/DATA2_1 , \U615/DATA2_2 , \U615/DATA2_3 ,
         \U615/DATA2_4 , \U615/DATA2_5 , \U615/DATA2_6 , \U615/DATA2_7 ,
         \U615/DATA2_8 , \U615/DATA2_9 , \U615/DATA2_10 , \U615/DATA2_11 ,
         \U615/DATA1_0 , \U615/DATA1_1 , \U615/DATA1_2 , \U615/DATA1_3 ,
         \U615/DATA1_4 , \U615/DATA1_5 , \U615/DATA1_6 , \U615/DATA1_7 ,
         \U615/DATA1_8 , \U615/DATA1_9 , \U615/DATA1_10 , \U615/DATA1_11 ,
         \U611/DATA1_0 , \U611/DATA1_1 , \U611/DATA1_2 , \U611/DATA1_3 ,
         \U611/DATA1_4 , \U611/DATA1_5 , \U611/DATA1_6 , \U611/DATA1_7 ,
         \U611/DATA1_8 , \U611/DATA1_9 , \U611/DATA1_10 , \U611/DATA1_11 ,
         \U610/DATA1_0 , \U610/DATA1_1 , \U610/DATA1_2 , \U610/DATA1_3 ,
         \U610/DATA1_4 , \U610/DATA1_5 , \U610/DATA1_6 , \U610/DATA1_7 ,
         \U610/DATA1_8 , \U610/DATA1_9 , \U610/DATA1_10 , \U610/DATA1_11 ,
         \U606/DATA1_0 , \U606/DATA1_1 , \U606/DATA1_2 , \U606/DATA1_3 ,
         \U606/DATA1_4 , \U606/DATA1_5 , \U606/DATA1_6 , \U606/DATA1_7 ,
         \U606/DATA1_8 , \U606/DATA1_9 , \U606/DATA1_10 , \U606/DATA1_11 ,
         \U605/DATA1_0 , \U605/DATA1_1 , \U605/DATA1_2 , \U605/DATA1_3 ,
         \U605/DATA1_4 , \U605/DATA1_5 , \U605/DATA1_6 , \U605/DATA1_7 ,
         \U605/DATA1_8 , \U605/DATA1_9 , \U605/DATA1_10 , \U605/DATA1_11 ,
         \U601/DATA1_0 , \U601/DATA1_1 , \U601/DATA1_2 , \U601/DATA1_3 ,
         \U601/DATA1_4 , \U601/DATA1_5 , \U601/DATA1_6 , \U601/DATA1_7 ,
         \U601/DATA1_8 , \U601/DATA1_9 , \U601/DATA1_10 , \U601/DATA1_11 ,
         \U600/DATA1_0 , \U600/DATA1_1 , \U600/DATA1_2 , \U600/DATA1_3 ,
         \U600/DATA1_4 , \U600/DATA1_5 , \U600/DATA1_6 , \U600/DATA1_7 ,
         \U600/DATA1_8 , \U600/DATA1_9 , \U600/DATA1_10 , \U600/DATA1_11 ,
         \U596/DATA1_0 , \U596/DATA1_1 , \U596/DATA1_2 , \U596/DATA1_3 ,
         \U596/DATA1_4 , \U596/DATA1_5 , \U596/DATA1_6 , \U596/DATA1_7 ,
         \U596/DATA1_8 , \U596/DATA1_9 , \U596/DATA1_10 , \U596/DATA1_11 ,
         \U595/DATA1_0 , \U595/DATA1_1 , \U595/DATA1_2 , \U595/DATA1_3 ,
         \U595/DATA1_4 , \U595/DATA1_5 , \U595/DATA1_6 , \U595/DATA1_7 ,
         \U595/DATA1_8 , \U595/DATA1_9 , \U595/DATA1_10 , \U595/DATA1_11 ,
         \U591/DATA1_0 , \U591/DATA1_1 , \U591/DATA1_2 , \U591/DATA1_3 ,
         \U591/DATA1_4 , \U591/DATA1_5 , \U591/DATA1_6 , \U591/DATA1_7 ,
         \U591/DATA1_8 , \U591/DATA1_9 , \U591/DATA1_10 , \U591/DATA1_11 ,
         \U590/DATA1_0 , \U590/DATA1_1 , \U590/DATA1_2 , \U590/DATA1_3 ,
         \U590/DATA1_4 , \U590/DATA1_5 , \U590/DATA1_6 , \U590/DATA1_7 ,
         \U590/DATA1_8 , \U590/DATA1_9 , \U590/DATA1_10 , \U590/DATA1_11 ,
         \U586/DATA1_0 , \U586/DATA1_1 , \U586/DATA1_2 , \U586/DATA1_3 ,
         \U586/DATA1_4 , \U586/DATA1_5 , \U586/DATA1_6 , \U586/DATA1_7 ,
         \U586/DATA1_8 , \U586/DATA1_9 , \U586/DATA1_10 , \U586/DATA1_11 ,
         \U585/DATA1_0 , \U585/DATA1_1 , \U585/DATA1_2 , \U585/DATA1_3 ,
         \U585/DATA1_4 , \U585/DATA1_5 , \U585/DATA1_6 , \U585/DATA1_7 ,
         \U585/DATA1_8 , \U585/DATA1_9 , \U585/DATA1_10 , \U585/DATA1_11 ,
         \U581/DATA1_0 , \U581/DATA1_1 , \U581/DATA1_2 , \U581/DATA1_3 ,
         \U581/DATA1_4 , \U581/DATA1_5 , \U581/DATA1_6 , \U581/DATA1_7 ,
         \U581/DATA1_8 , \U581/DATA1_9 , \U581/DATA1_10 , \U581/DATA1_11 ,
         \U580/DATA1_0 , \U580/DATA1_1 , \U580/DATA1_2 , \U580/DATA1_3 ,
         \U580/DATA1_4 , \U580/DATA1_5 , \U580/DATA1_6 , \U580/DATA1_7 ,
         \U580/DATA1_8 , \U580/DATA1_9 , \U580/DATA1_10 , \U580/DATA1_11 ,
         \U576/DATA1_0 , \U576/DATA1_1 , \U576/DATA1_2 , \U576/DATA1_3 ,
         \U576/DATA1_4 , \U576/DATA1_5 , \U576/DATA1_6 , \U576/DATA1_7 ,
         \U576/DATA1_8 , \U576/DATA1_9 , \U576/DATA1_10 , \U576/DATA1_11 ,
         \U575/DATA1_0 , \U575/DATA1_1 , \U575/DATA1_2 , \U575/DATA1_3 ,
         \U575/DATA1_4 , \U575/DATA1_5 , \U575/DATA1_6 , \U575/DATA1_7 ,
         \U575/DATA1_8 , \U575/DATA1_9 , \U575/DATA1_10 , \U575/DATA1_11 ,
         \U571/DATA1_0 , \U571/DATA1_1 , \U571/DATA1_2 , \U571/DATA1_3 ,
         \U571/DATA1_4 , \U571/DATA1_5 , \U571/DATA1_6 , \U571/DATA1_7 ,
         \U571/DATA1_8 , \U571/DATA1_9 , \U571/DATA1_10 , \U571/DATA1_11 ,
         \U570/DATA1_0 , \U570/DATA1_1 , \U570/DATA1_2 , \U570/DATA1_3 ,
         \U570/DATA1_4 , \U570/DATA1_5 , \U570/DATA1_6 , \U570/DATA1_7 ,
         \U570/DATA1_8 , \U570/DATA1_9 , \U570/DATA1_10 , \U570/DATA1_11 ,
         \U565/DATA2_0 , \U565/DATA2_1 , \U565/DATA2_2 , \U565/DATA2_3 ,
         \U565/DATA2_4 , \U565/DATA2_5 , \U565/DATA2_6 , \U565/DATA2_7 ,
         \U565/DATA2_8 , \U565/DATA2_9 , \U565/DATA1_0 , \U565/DATA1_1 ,
         \U565/DATA1_2 , \U565/DATA1_3 , \U565/DATA1_4 , \U565/DATA1_5 ,
         \U565/DATA1_6 , \U565/DATA1_7 , \U565/DATA1_8 , \U565/DATA1_9 ,
         \U565/DATA1_10 , \U565/DATA1_11 , \U553/DATA2_0 , \U553/DATA2_1 ,
         \U553/DATA2_2 , \U553/DATA2_3 , \U553/DATA2_4 , \U553/DATA2_5 ,
         \U553/DATA2_6 , \U553/DATA2_7 , \U553/DATA2_8 , \U553/DATA2_9 ,
         \U553/DATA2_10 , \U553/DATA2_11 , \U553/DATA1_0 , \U553/DATA1_1 ,
         \U553/DATA1_2 , \U553/DATA1_3 , \U553/DATA1_4 , \U553/DATA1_5 ,
         \U553/DATA1_6 , \U553/DATA1_7 , \U553/DATA1_8 , \U553/DATA1_9 ,
         \U553/DATA1_10 , \U553/DATA1_11 , \U548/DATA1_0 , \U548/DATA1_1 ,
         \U548/DATA1_2 , \U548/DATA1_3 , \U548/DATA1_4 , \U548/DATA1_5 ,
         \U548/DATA1_6 , \U548/DATA1_7 , \U548/DATA1_8 , \U548/DATA1_9 ,
         \U548/DATA1_10 , \U548/DATA1_11 , \U543/DATA1_0 , \U543/DATA1_1 ,
         \U543/DATA1_2 , \U543/DATA1_3 , \U543/DATA1_4 , \U543/DATA1_5 ,
         \U543/DATA1_6 , \U543/DATA1_7 , \U543/DATA1_8 , \U543/DATA1_9 ,
         \U543/DATA1_10 , \U543/DATA1_11 , \U538/DATA1_0 , \U538/DATA1_1 ,
         \U538/DATA1_2 , \U538/DATA1_3 , \U538/DATA1_4 , \U538/DATA1_5 ,
         \U538/DATA1_6 , \U538/DATA1_7 , \U538/DATA1_8 , \U538/DATA1_9 ,
         \U538/DATA1_10 , \U538/DATA1_11 , \U533/DATA1_0 , \U533/DATA1_1 ,
         \U533/DATA1_2 , \U533/DATA1_3 , \U533/DATA1_4 , \U533/DATA1_5 ,
         \U533/DATA1_6 , \U533/DATA1_7 , \U533/DATA1_8 , \U533/DATA1_9 ,
         \U533/DATA1_10 , \U533/DATA1_11 , \U528/DATA1_0 , \U528/DATA1_1 ,
         \U528/DATA1_2 , \U528/DATA1_3 , \U528/DATA1_4 , \U528/DATA1_5 ,
         \U528/DATA1_6 , \U528/DATA1_7 , \U528/DATA1_8 , \U528/DATA1_9 ,
         \U528/DATA1_10 , \U528/DATA1_11 , \U523/DATA1_0 , \U523/DATA1_1 ,
         \U523/DATA1_2 , \U523/DATA1_3 , \U523/DATA1_4 , \U523/DATA1_5 ,
         \U523/DATA1_6 , \U523/DATA1_7 , \U523/DATA1_8 , \U523/DATA1_9 ,
         \U523/DATA1_10 , \U523/DATA1_11 , \U518/DATA1_0 , \U518/DATA1_1 ,
         \U518/DATA1_2 , \U518/DATA1_3 , \U518/DATA1_4 , \U518/DATA1_5 ,
         \U518/DATA1_6 , \U518/DATA1_7 , \U518/DATA1_8 , \U518/DATA1_9 ,
         \U518/DATA1_10 , \U518/DATA1_11 , \U513/DATA1_0 , \U513/DATA1_1 ,
         \U513/DATA1_2 , \U513/DATA1_3 , \U513/DATA1_4 , \U513/DATA1_5 ,
         \U513/DATA1_6 , \U513/DATA1_7 , \U513/DATA1_8 , \U513/DATA1_9 ,
         \U513/DATA1_10 , \U513/DATA1_11 , \U508/DATA1_0 , \U508/DATA1_1 ,
         \U508/DATA1_2 , \U508/DATA1_3 , \U508/DATA1_4 , \U508/DATA1_5 ,
         \U508/DATA1_6 , \U508/DATA1_7 , \U508/DATA1_8 , \U508/DATA1_9 ,
         \U508/DATA1_10 , \U508/DATA1_11 , \U503/DATA2_0 , \U503/DATA2_1 ,
         \U503/DATA2_2 , \U503/DATA2_3 , \U503/DATA2_4 , \U503/DATA2_5 ,
         \U503/DATA2_6 , \U503/DATA2_7 , \U503/DATA2_8 , \U503/DATA2_9 ,
         \U503/DATA1_0 , \U503/DATA1_1 , \U503/DATA1_2 , \U503/DATA1_3 ,
         \U503/DATA1_4 , \U503/DATA1_5 , \U503/DATA1_6 , \U503/DATA1_7 ,
         \U503/DATA1_8 , \U503/DATA1_9 , \U503/DATA1_10 , \U503/DATA1_11 ,
         \U500/DATA2_0 , \U500/DATA2_1 , \U500/DATA2_2 , \U500/DATA2_3 ,
         \U500/DATA2_4 , \U500/DATA2_5 , \U500/DATA2_6 , \U500/DATA2_7 ,
         \U500/DATA2_8 , \U500/DATA2_9 , \U500/DATA2_10 , \U500/DATA2_11 ,
         \U500/DATA1_0 , \U500/DATA1_1 , \U500/DATA1_2 , \U500/DATA1_3 ,
         \U500/DATA1_4 , \U500/DATA1_5 , \U500/DATA1_6 , \U500/DATA1_7 ,
         \U500/DATA1_8 , \U500/DATA1_9 , \U500/DATA1_10 , \U500/DATA1_11 ,
         \U495/DATA1_0 , \U495/DATA1_1 , \U495/DATA1_2 , \U495/DATA1_3 ,
         \U495/DATA1_4 , \U495/DATA1_5 , \U495/DATA1_6 , \U495/DATA1_7 ,
         \U495/DATA1_8 , \U495/DATA1_9 , \U495/DATA1_10 , \U495/DATA1_11 ,
         \U490/DATA1_0 , \U490/DATA1_1 , \U490/DATA1_2 , \U490/DATA1_3 ,
         \U490/DATA1_4 , \U490/DATA1_5 , \U490/DATA1_6 , \U490/DATA1_7 ,
         \U490/DATA1_8 , \U490/DATA1_9 , \U490/DATA1_10 , \U490/DATA1_11 ,
         \U485/DATA1_0 , \U485/DATA1_1 , \U485/DATA1_2 , \U485/DATA1_3 ,
         \U485/DATA1_4 , \U485/DATA1_5 , \U485/DATA1_6 , \U485/DATA1_7 ,
         \U485/DATA1_8 , \U485/DATA1_9 , \U485/DATA1_10 , \U485/DATA1_11 ,
         \U480/DATA1_0 , \U480/DATA1_1 , \U480/DATA1_2 , \U480/DATA1_3 ,
         \U480/DATA1_4 , \U480/DATA1_5 , \U480/DATA1_6 , \U480/DATA1_7 ,
         \U480/DATA1_8 , \U480/DATA1_9 , \U480/DATA1_10 , \U480/DATA1_11 ,
         \U475/DATA1_0 , \U475/DATA1_1 , \U475/DATA1_2 , \U475/DATA1_3 ,
         \U475/DATA1_4 , \U475/DATA1_5 , \U475/DATA1_6 , \U475/DATA1_7 ,
         \U475/DATA1_8 , \U475/DATA1_9 , \U475/DATA1_10 , \U475/DATA1_11 ,
         \U470/DATA1_0 , \U470/DATA1_1 , \U470/DATA1_2 , \U470/DATA1_3 ,
         \U470/DATA1_4 , \U470/DATA1_5 , \U470/DATA1_6 , \U470/DATA1_7 ,
         \U470/DATA1_8 , \U470/DATA1_9 , \U470/DATA1_10 , \U470/DATA1_11 ,
         \U465/DATA1_0 , \U465/DATA1_1 , \U465/DATA1_2 , \U465/DATA1_3 ,
         \U465/DATA1_4 , \U465/DATA1_5 , \U465/DATA1_6 , \U465/DATA1_7 ,
         \U465/DATA1_8 , \U465/DATA1_9 , \U465/DATA1_10 , \U465/DATA1_11 ,
         \U460/DATA1_0 , \U460/DATA1_1 , \U460/DATA1_2 , \U460/DATA1_3 ,
         \U460/DATA1_4 , \U460/DATA1_5 , \U460/DATA1_6 , \U460/DATA1_7 ,
         \U460/DATA1_8 , \U460/DATA1_9 , \U460/DATA1_10 , \U460/DATA1_11 ,
         \U455/DATA1_0 , \U455/DATA1_1 , \U455/DATA1_2 , \U455/DATA1_3 ,
         \U455/DATA1_4 , \U455/DATA1_5 , \U455/DATA1_6 , \U455/DATA1_7 ,
         \U455/DATA1_8 , \U455/DATA1_9 , \U455/DATA1_10 , \U455/DATA1_11 ,
         \U450/DATA2_0 , \U450/DATA2_1 , \U450/DATA2_2 , \U450/DATA2_3 ,
         \U450/DATA2_4 , \U450/DATA2_5 , \U450/DATA2_6 , \U450/DATA2_7 ,
         \U450/DATA2_8 , \U450/DATA2_9 , \U450/DATA1_0 , \U450/DATA1_1 ,
         \U450/DATA1_2 , \U450/DATA1_3 , \U450/DATA1_4 , \U450/DATA1_5 ,
         \U450/DATA1_6 , \U450/DATA1_7 , \U450/DATA1_8 , \U450/DATA1_9 ,
         \U450/DATA1_10 , \U450/DATA1_11 , \U444/DATA2_0 , \U444/DATA2_1 ,
         \U444/DATA2_2 , \U444/DATA2_3 , \U444/DATA2_4 , \U444/DATA2_5 ,
         \U444/DATA2_6 , \U444/DATA2_7 , \U444/DATA2_8 , \U444/DATA2_9 ,
         \U444/DATA2_10 , \U444/DATA2_11 , \U444/DATA1_0 , \U444/DATA1_1 ,
         \U444/DATA1_2 , \U444/DATA1_3 , \U444/DATA1_4 , \U444/DATA1_5 ,
         \U444/DATA1_6 , \U444/DATA1_7 , \U444/DATA1_8 , \U444/DATA1_9 ,
         \U444/DATA1_10 , \U444/DATA1_11 , \U439/DATA1_0 , \U439/DATA1_1 ,
         \U439/DATA1_2 , \U439/DATA1_3 , \U439/DATA1_4 , \U439/DATA1_5 ,
         \U439/DATA1_6 , \U439/DATA1_7 , \U439/DATA1_8 , \U439/DATA1_9 ,
         \U439/DATA1_10 , \U439/DATA1_11 , \U434/DATA1_0 , \U434/DATA1_1 ,
         \U434/DATA1_2 , \U434/DATA1_3 , \U434/DATA1_4 , \U434/DATA1_5 ,
         \U434/DATA1_6 , \U434/DATA1_7 , \U434/DATA1_8 , \U434/DATA1_9 ,
         \U434/DATA1_10 , \U434/DATA1_11 , \U429/DATA1_0 , \U429/DATA1_1 ,
         \U429/DATA1_2 , \U429/DATA1_3 , \U429/DATA1_4 , \U429/DATA1_5 ,
         \U429/DATA1_6 , \U429/DATA1_7 , \U429/DATA1_8 , \U429/DATA1_9 ,
         \U429/DATA1_10 , \U429/DATA1_11 , \U424/DATA1_0 , \U424/DATA1_1 ,
         \U424/DATA1_2 , \U424/DATA1_3 , \U424/DATA1_4 , \U424/DATA1_5 ,
         \U424/DATA1_6 , \U424/DATA1_7 , \U424/DATA1_8 , \U424/DATA1_9 ,
         \U424/DATA1_10 , \U424/DATA1_11 , \U419/DATA1_0 , \U419/DATA1_1 ,
         \U419/DATA1_2 , \U419/DATA1_3 , \U419/DATA1_4 , \U419/DATA1_5 ,
         \U419/DATA1_6 , \U419/DATA1_7 , \U419/DATA1_8 , \U419/DATA1_9 ,
         \U419/DATA1_10 , \U419/DATA1_11 , \U414/DATA1_0 , \U414/DATA1_1 ,
         \U414/DATA1_2 , \U414/DATA1_3 , \U414/DATA1_4 , \U414/DATA1_5 ,
         \U414/DATA1_6 , \U414/DATA1_7 , \U414/DATA1_8 , \U414/DATA1_9 ,
         \U414/DATA1_10 , \U414/DATA1_11 , \U409/DATA1_0 , \U409/DATA1_1 ,
         \U409/DATA1_2 , \U409/DATA1_3 , \U409/DATA1_4 , \U409/DATA1_5 ,
         \U409/DATA1_6 , \U409/DATA1_7 , \U409/DATA1_8 , \U409/DATA1_9 ,
         \U409/DATA1_10 , \U409/DATA1_11 , \U404/DATA1_0 , \U404/DATA1_1 ,
         \U404/DATA1_2 , \U404/DATA1_3 , \U404/DATA1_4 , \U404/DATA1_5 ,
         \U404/DATA1_6 , \U404/DATA1_7 , \U404/DATA1_8 , \U404/DATA1_9 ,
         \U404/DATA1_10 , \U404/DATA1_11 , \U399/DATA1_0 , \U399/DATA1_1 ,
         \U399/DATA1_2 , \U399/DATA1_3 , \U399/DATA1_4 , \U399/DATA1_5 ,
         \U399/DATA1_6 , \U399/DATA1_7 , \U399/DATA1_8 , \U399/DATA1_9 ,
         \U399/DATA1_10 , \U399/DATA1_11 , \U394/DATA2_0 , \U394/DATA2_1 ,
         \U394/DATA2_2 , \U394/DATA2_3 , \U394/DATA2_4 , \U394/DATA2_5 ,
         \U394/DATA2_6 , \U394/DATA2_7 , \U394/DATA2_8 , \U394/DATA2_9 ,
         \U394/DATA1_0 , \U394/DATA1_1 , \U394/DATA1_2 , \U394/DATA1_3 ,
         \U394/DATA1_4 , \U394/DATA1_5 , \U394/DATA1_6 , \U394/DATA1_7 ,
         \U394/DATA1_8 , \U394/DATA1_9 , \U394/DATA1_10 , \U394/DATA1_11 ,
         \U391/DATA2_0 , \U391/DATA2_1 , \U391/DATA2_2 , \U391/DATA2_3 ,
         \U391/DATA2_4 , \U391/DATA2_5 , \U391/DATA2_6 , \U391/DATA2_7 ,
         \U391/DATA2_8 , \U391/DATA2_9 , \U391/DATA2_10 , \U391/DATA2_11 ,
         \U391/DATA1_0 , \U391/DATA1_1 , \U391/DATA1_2 , \U391/DATA1_3 ,
         \U391/DATA1_4 , \U391/DATA1_5 , \U391/DATA1_6 , \U391/DATA1_7 ,
         \U391/DATA1_8 , \U391/DATA1_9 , \U391/DATA1_10 , \U391/DATA1_11 ,
         \U386/DATA1_0 , \U386/DATA1_1 , \U386/DATA1_2 , \U386/DATA1_3 ,
         \U386/DATA1_4 , \U386/DATA1_5 , \U386/DATA1_6 , \U386/DATA1_7 ,
         \U386/DATA1_8 , \U386/DATA1_9 , \U386/DATA1_10 , \U386/DATA1_11 ,
         \U381/DATA1_0 , \U381/DATA1_1 , \U381/DATA1_2 , \U381/DATA1_3 ,
         \U381/DATA1_4 , \U381/DATA1_5 , \U381/DATA1_6 , \U381/DATA1_7 ,
         \U381/DATA1_8 , \U381/DATA1_9 , \U381/DATA1_10 , \U381/DATA1_11 ,
         \U376/DATA1_0 , \U376/DATA1_1 , \U376/DATA1_2 , \U376/DATA1_3 ,
         \U376/DATA1_4 , \U376/DATA1_5 , \U376/DATA1_6 , \U376/DATA1_7 ,
         \U376/DATA1_8 , \U376/DATA1_9 , \U376/DATA1_10 , \U376/DATA1_11 ,
         \U371/DATA1_0 , \U371/DATA1_1 , \U371/DATA1_2 , \U371/DATA1_3 ,
         \U371/DATA1_4 , \U371/DATA1_5 , \U371/DATA1_6 , \U371/DATA1_7 ,
         \U371/DATA1_8 , \U371/DATA1_9 , \U371/DATA1_10 , \U371/DATA1_11 ,
         \U366/DATA1_0 , \U366/DATA1_1 , \U366/DATA1_2 , \U366/DATA1_3 ,
         \U366/DATA1_4 , \U366/DATA1_5 , \U366/DATA1_6 , \U366/DATA1_7 ,
         \U366/DATA1_8 , \U366/DATA1_9 , \U366/DATA1_10 , \U366/DATA1_11 ,
         \U361/DATA1_3 , \U361/DATA1_4 , \U361/DATA1_5 , \U361/DATA1_6 ,
         \U361/DATA1_7 , \U361/DATA1_8 , \U361/DATA1_9 , \U361/DATA1_10 ,
         \U361/DATA1_11 , \U356/DATA1_1 , \U356/DATA1_2 , \U356/DATA1_3 ,
         \U356/DATA1_4 , \U356/DATA1_5 , \U356/DATA1_6 , \U356/DATA1_7 ,
         \U356/DATA1_8 , \U356/DATA1_9 , \U356/DATA1_10 , \U356/DATA1_11 ,
         \U351/DATA1_1 , \U351/DATA1_2 , \U351/DATA1_3 , \U351/DATA1_4 ,
         \U351/DATA1_5 , \U351/DATA1_6 , \U351/DATA1_7 , \U351/DATA1_8 ,
         \U351/DATA1_9 , \U351/DATA1_10 , \U351/DATA1_11 , \U346/DATA1_5 ,
         \U346/DATA1_6 , \U346/DATA1_7 , \U346/DATA1_8 , \U346/DATA1_9 ,
         \U346/DATA1_10 , \U346/DATA1_11 , \U341/DATA2_1 , \U341/DATA2_2 ,
         \U341/DATA2_3 , \U341/DATA2_4 , \U341/DATA2_5 , \U341/DATA2_6 ,
         \U341/DATA2_7 , \U341/DATA2_8 , \U341/DATA2_9 , \U341/DATA1_1 ,
         \U341/DATA1_2 , \U341/DATA1_3 , \U341/DATA1_4 , \U341/DATA1_5 ,
         \U341/DATA1_6 , \U341/DATA1_7 , \U341/DATA1_8 , \U341/DATA1_9 ,
         \U341/DATA1_10 , \U341/DATA1_11 , \U332/DATA2_1 , \U332/DATA2_2 ,
         \U332/DATA2_3 , \U332/DATA2_4 , \U332/DATA2_5 , \U332/DATA2_6 ,
         \U332/DATA2_7 , \U332/DATA2_8 , \U332/DATA2_9 , \U332/DATA2_10 ,
         \U332/DATA2_11 , \U332/DATA1_1 , \U332/DATA1_2 , \U332/DATA1_3 ,
         \U332/DATA1_4 , \U332/DATA1_5 , \U332/DATA1_6 , \U332/DATA1_7 ,
         \U332/DATA1_8 , \U332/DATA1_9 , \U332/DATA1_10 , \U332/DATA1_11 ,
         \U327/DATA1_2 , \U327/DATA1_3 , \U327/DATA1_4 , \U327/DATA1_5 ,
         \U327/DATA1_6 , \U327/DATA1_7 , \U327/DATA1_8 , \U327/DATA1_9 ,
         \U327/DATA1_10 , \U327/DATA1_11 , \U322/DATA1_3 , \U322/DATA1_4 ,
         \U322/DATA1_5 , \U322/DATA1_6 , \U322/DATA1_7 , \U322/DATA1_8 ,
         \U322/DATA1_9 , \U322/DATA1_10 , \U322/DATA1_11 , \U317/DATA1_1 ,
         \U317/DATA1_2 , \U317/DATA1_3 , \U317/DATA1_4 , \U317/DATA1_5 ,
         \U317/DATA1_6 , \U317/DATA1_7 , \U317/DATA1_8 , \U317/DATA1_9 ,
         \U317/DATA1_10 , \U317/DATA1_11 , \U312/DATA1_1 , \U312/DATA1_2 ,
         \U312/DATA1_3 , \U312/DATA1_4 , \U312/DATA1_5 , \U312/DATA1_6 ,
         \U312/DATA1_7 , \U312/DATA1_8 , \U312/DATA1_9 , \U312/DATA1_10 ,
         \U312/DATA1_11 , \U307/DATA1_5 , \U307/DATA1_6 , \U307/DATA1_7 ,
         \U307/DATA1_8 , \U307/DATA1_9 , \U307/DATA1_10 , \U307/DATA1_11 ,
         \U302/DATA1_1 , \U302/DATA1_2 , \U302/DATA1_3 , \U302/DATA1_4 ,
         \U302/DATA1_5 , \U302/DATA1_6 , \U302/DATA1_7 , \U302/DATA1_8 ,
         \U302/DATA1_9 , \U302/DATA1_10 , \U302/DATA1_11 , \U297/DATA1_7 ,
         \U297/DATA1_8 , \U297/DATA1_9 , \U297/DATA1_10 , \U297/DATA1_11 ,
         \U292/DATA1_1 , \U292/DATA1_2 , \U292/DATA1_3 , \U292/DATA1_4 ,
         \U292/DATA1_5 , \U292/DATA1_6 , \U292/DATA1_7 , \U292/DATA1_8 ,
         \U292/DATA1_9 , \U292/DATA1_10 , \U292/DATA1_11 , \U287/DATA1_2 ,
         \U287/DATA1_3 , \U287/DATA1_4 , \U287/DATA1_5 , \U287/DATA1_6 ,
         \U287/DATA1_7 , \U287/DATA1_8 , \U287/DATA1_9 , \U287/DATA1_10 ,
         \U287/DATA1_11 , \U282/DATA2_1 , \U282/DATA2_2 , \U282/DATA2_3 ,
         \U282/DATA2_4 , \U282/DATA2_5 , \U282/DATA2_6 , \U282/DATA2_7 ,
         \U282/DATA2_8 , \U282/DATA2_9 , \U282/DATA1_1 , \U282/DATA1_2 ,
         \U282/DATA1_3 , \U282/DATA1_4 , \U282/DATA1_5 , \U282/DATA1_6 ,
         \U282/DATA1_7 , \U282/DATA1_8 , \U282/DATA1_9 , \U282/DATA1_10 ,
         \U282/DATA1_11 , \U279/DATA2_1 , \U279/DATA2_2 , \U279/DATA2_3 ,
         \U279/DATA2_4 , \U279/DATA2_5 , \U279/DATA2_6 , \U279/DATA2_7 ,
         \U279/DATA2_8 , \U279/DATA2_9 , \U279/DATA2_10 , \U279/DATA2_11 ,
         \U279/DATA1_1 , \U279/DATA1_2 , \U279/DATA1_3 , \U279/DATA1_4 ,
         \U279/DATA1_5 , \U279/DATA1_6 , \U279/DATA1_7 , \U279/DATA1_8 ,
         \U279/DATA1_9 , \U279/DATA1_10 , \U279/DATA1_11 , \U274/DATA1_2 ,
         \U274/DATA1_3 , \U274/DATA1_4 , \U274/DATA1_5 , \U274/DATA1_6 ,
         \U274/DATA1_7 , \U274/DATA1_8 , \U274/DATA1_9 , \U274/DATA1_10 ,
         \U274/DATA1_11 , \U269/DATA1_1 , \U269/DATA1_2 , \U269/DATA1_3 ,
         \U269/DATA1_4 , \U269/DATA1_5 , \U269/DATA1_6 , \U269/DATA1_7 ,
         \U269/DATA1_8 , \U269/DATA1_9 , \U269/DATA1_10 , \U269/DATA1_11 ,
         \U264/DATA1_1 , \U264/DATA1_2 , \U264/DATA1_3 , \U264/DATA1_4 ,
         \U264/DATA1_5 , \U264/DATA1_6 , \U264/DATA1_7 , \U264/DATA1_8 ,
         \U264/DATA1_9 , \U264/DATA1_10 , \U264/DATA1_11 , \U254/DATA1_1 ,
         \U254/DATA1_2 , \U254/DATA1_3 , \U254/DATA1_4 , \U254/DATA1_5 ,
         \U254/DATA1_6 , \U254/DATA1_7 , \U254/DATA1_8 , \U254/DATA1_9 ,
         \U254/DATA1_10 , \U254/DATA1_11 , \U249/DATA1_2 , \U249/DATA1_3 ,
         \U249/DATA1_4 , \U249/DATA1_5 , \U249/DATA1_6 , \U249/DATA1_7 ,
         \U249/DATA1_8 , \U249/DATA1_9 , \U249/DATA1_10 , \U249/DATA1_11 ,
         \U244/DATA1_3 , \U244/DATA1_4 , \U244/DATA1_5 , \U244/DATA1_6 ,
         \U244/DATA1_7 , \U244/DATA1_8 , \U244/DATA1_9 , \U244/DATA1_10 ,
         \U244/DATA1_11 , \U239/DATA1_1 , \U239/DATA1_2 , \U239/DATA1_3 ,
         \U239/DATA1_4 , \U239/DATA1_5 , \U239/DATA1_6 , \U239/DATA1_7 ,
         \U239/DATA1_8 , \U239/DATA1_9 , \U239/DATA1_10 , \U239/DATA1_11 ,
         \U234/DATA1_1 , \U234/DATA1_2 , \U234/DATA1_3 , \U234/DATA1_4 ,
         \U234/DATA1_5 , \U234/DATA1_6 , \U234/DATA1_7 , \U234/DATA1_8 ,
         \U234/DATA1_9 , \U234/DATA1_10 , \U234/DATA1_11 , \U229/DATA2_6 ,
         \U229/DATA2_7 , \U229/DATA2_8 , \U229/DATA2_9 , \U229/DATA1_6 ,
         \U229/DATA1_7 , \U229/DATA1_8 , \U229/DATA1_9 , \U229/DATA1_10 ,
         \U229/DATA1_11 , \U223/DATA2_6 , \U223/DATA2_7 , \U223/DATA2_8 ,
         \U223/DATA2_9 , \U223/DATA2_10 , \U223/DATA2_11 , \U223/DATA1_6 ,
         \U223/DATA1_7 , \U223/DATA1_8 , \U223/DATA1_9 , \U223/DATA1_10 ,
         \U223/DATA1_11 , \U218/DATA1_6 , \U218/DATA1_7 , \U218/DATA1_8 ,
         \U218/DATA1_9 , \U218/DATA1_10 , \U218/DATA1_11 , \U213/DATA1_6 ,
         \U213/DATA1_7 , \U213/DATA1_8 , \U213/DATA1_9 , \U213/DATA1_10 ,
         \U213/DATA1_11 , \U208/DATA1_6 , \U208/DATA1_7 , \U208/DATA1_8 ,
         \U208/DATA1_9 , \U208/DATA1_10 , \U208/DATA1_11 , \U203/DATA1_7 ,
         \U203/DATA1_8 , \U203/DATA1_9 , \U203/DATA1_10 , \U203/DATA1_11 ,
         \U198/DATA1_7 , \U198/DATA1_8 , \U198/DATA1_9 , \U198/DATA1_10 ,
         \U198/DATA1_11 , \U193/DATA1_7 , \U193/DATA1_8 , \U193/DATA1_9 ,
         \U193/DATA1_10 , \U193/DATA1_11 , \U188/DATA1_7 , \U188/DATA1_8 ,
         \U188/DATA1_9 , \U188/DATA1_10 , \U188/DATA1_11 , \U183/DATA1_7 ,
         \U183/DATA1_8 , \U183/DATA1_9 , \U183/DATA1_10 , \U183/DATA1_11 ,
         \U178/DATA1_7 , \U178/DATA1_8 , \U178/DATA1_9 , \U178/DATA1_10 ,
         \U178/DATA1_11 , \U173/DATA2_2 , \U173/DATA2_3 , \U173/DATA2_4 ,
         \U173/DATA2_5 , \U173/DATA2_6 , \U173/DATA2_7 , \U173/DATA2_8 ,
         \U173/DATA2_9 , \U173/DATA1_2 , \U173/DATA1_3 , \U173/DATA1_4 ,
         \U173/DATA1_5 , \U173/DATA1_6 , \U173/DATA1_7 , \U173/DATA1_8 ,
         \U173/DATA1_9 , \U173/DATA1_10 , \U173/DATA1_11 , \U170/DATA2_2 ,
         \U170/DATA2_3 , \U170/DATA2_4 , \U170/DATA2_5 , \U170/DATA2_6 ,
         \U170/DATA2_7 , \U170/DATA2_8 , \U170/DATA2_9 , \U170/DATA2_10 ,
         \U170/DATA2_11 , \U170/DATA1_2 , \U170/DATA1_3 , \U170/DATA1_4 ,
         \U170/DATA1_5 , \U170/DATA1_6 , \U170/DATA1_7 , \U170/DATA1_8 ,
         \U170/DATA1_9 , \U170/DATA1_10 , \U170/DATA1_11 , \U165/DATA1_2 ,
         \U165/DATA1_3 , \U165/DATA1_4 , \U165/DATA1_5 , \U165/DATA1_6 ,
         \U165/DATA1_7 , \U165/DATA1_8 , \U165/DATA1_9 , \U165/DATA1_10 ,
         \U165/DATA1_11 , \U160/DATA1_2 , \U160/DATA1_3 , \U160/DATA1_4 ,
         \U160/DATA1_5 , \U160/DATA1_6 , \U160/DATA1_7 , \U160/DATA1_8 ,
         \U160/DATA1_9 , \U160/DATA1_10 , \U160/DATA1_11 , \U155/DATA1_2 ,
         \U155/DATA1_3 , \U155/DATA1_4 , \U155/DATA1_5 , \U155/DATA1_6 ,
         \U155/DATA1_7 , \U155/DATA1_8 , \U155/DATA1_9 , \U155/DATA1_10 ,
         \U155/DATA1_11 , \U150/DATA1_2 , \U150/DATA1_3 , \U150/DATA1_4 ,
         \U150/DATA1_5 , \U150/DATA1_6 , \U150/DATA1_7 , \U150/DATA1_8 ,
         \U150/DATA1_9 , \U150/DATA1_10 , \U150/DATA1_11 , \U145/DATA1_2 ,
         \U145/DATA1_3 , \U145/DATA1_4 , \U145/DATA1_5 , \U145/DATA1_6 ,
         \U145/DATA1_7 , \U145/DATA1_8 , \U145/DATA1_9 , \U145/DATA1_10 ,
         \U145/DATA1_11 , \U140/DATA1_0 , \U140/DATA1_1 , \U140/DATA1_2 ,
         \U140/DATA1_3 , \U140/DATA1_4 , \U140/DATA1_5 , \U140/DATA1_6 ,
         \U140/DATA1_7 , \U140/DATA1_8 , \U140/DATA1_9 , \U140/DATA1_10 ,
         \U140/DATA1_11 , \U135/DATA1_0 , \U135/DATA1_1 , \U135/DATA1_2 ,
         \U135/DATA1_3 , \U135/DATA1_4 , \U135/DATA1_5 , \U135/DATA1_6 ,
         \U135/DATA1_7 , \U135/DATA1_8 , \U135/DATA1_9 , \U135/DATA1_10 ,
         \U135/DATA1_11 , \U130/DATA1_0 , \U130/DATA1_1 , \U130/DATA1_2 ,
         \U130/DATA1_3 , \U130/DATA1_4 , \U130/DATA1_5 , \U130/DATA1_6 ,
         \U130/DATA1_7 , \U130/DATA1_8 , \U130/DATA1_9 , \U130/DATA1_10 ,
         \U130/DATA1_11 , \U125/DATA1_0 , \U125/DATA1_1 , \U125/DATA1_2 ,
         \U125/DATA1_3 , \U125/DATA1_4 , \U125/DATA1_5 , \U125/DATA1_6 ,
         \U125/DATA1_7 , \U125/DATA1_8 , \U125/DATA1_9 , \U125/DATA1_10 ,
         \U125/DATA1_11 , \U120/DATA2_0 , \U120/DATA2_1 , \U120/DATA2_2 ,
         \U120/DATA2_3 , \U120/DATA2_4 , \U120/DATA2_5 , \U120/DATA2_6 ,
         \U120/DATA2_7 , \U120/DATA2_8 , \U120/DATA1_0 , \U120/DATA1_1 ,
         \U120/DATA1_2 , \U120/DATA1_3 , \U120/DATA1_4 , \U120/DATA1_5 ,
         \U120/DATA1_6 , \U120/DATA1_7 , \U120/DATA1_8 , \U120/DATA1_9 ,
         \U120/DATA1_10 , \U120/DATA1_11 , \U108/DATA2_0 , \U108/DATA2_1 ,
         \U108/DATA2_2 , \U108/DATA2_3 , \U108/DATA2_4 , \U108/DATA2_5 ,
         \U108/DATA2_6 , \U108/DATA2_7 , \U108/DATA2_8 , \U108/DATA2_9 ,
         \U108/DATA2_10 , \U108/DATA2_11 , \U108/DATA1_0 , \U108/DATA1_1 ,
         \U108/DATA1_2 , \U108/DATA1_3 , \U108/DATA1_4 , \U108/DATA1_5 ,
         \U108/DATA1_6 , \U108/DATA1_7 , \U108/DATA1_8 , \U108/DATA1_9 ,
         \U108/DATA1_10 , \U108/DATA1_11 , \U103/DATA1_0 , \U103/DATA1_1 ,
         \U103/DATA1_2 , \U103/DATA1_3 , \U103/DATA1_4 , \U103/DATA1_5 ,
         \U103/DATA1_6 , \U103/DATA1_7 , \U103/DATA1_8 , \U103/DATA1_9 ,
         \U103/DATA1_10 , \U103/DATA1_11 , \U98/DATA1_0 , \U98/DATA1_1 ,
         \U98/DATA1_2 , \U98/DATA1_3 , \U98/DATA1_4 , \U98/DATA1_5 ,
         \U98/DATA1_6 , \U98/DATA1_7 , \U98/DATA1_8 , \U98/DATA1_9 ,
         \U98/DATA1_10 , \U98/DATA1_11 , \U93/DATA1_5 , \U93/DATA1_6 ,
         \U93/DATA1_7 , \U93/DATA1_8 , \U93/DATA1_9 , \U93/DATA1_10 ,
         \U93/DATA1_11 , \U88/DATA1_1 , \U88/DATA1_2 , \U88/DATA1_3 ,
         \U88/DATA1_4 , \U88/DATA1_5 , \U88/DATA1_6 , \U88/DATA1_7 ,
         \U88/DATA1_8 , \U88/DATA1_9 , \U88/DATA1_10 , \U88/DATA1_11 ,
         \U83/DATA1_4 , \U83/DATA1_5 , \U83/DATA1_6 , \U83/DATA1_7 ,
         \U83/DATA1_8 , \U83/DATA1_9 , \U83/DATA1_10 , \U83/DATA1_11 ,
         \U78/DATA1_9 , \U78/DATA1_10 , \U78/DATA1_11 , \U73/DATA1_1 ,
         \U73/DATA1_2 , \U73/DATA1_3 , \U73/DATA1_4 , \U73/DATA1_5 ,
         \U73/DATA1_6 , \U73/DATA1_7 , \U73/DATA1_8 , \U73/DATA1_9 ,
         \U73/DATA1_10 , \U73/DATA1_11 , \U68/DATA1_6 , \U68/DATA1_7 ,
         \U68/DATA1_8 , \U68/DATA1_9 , \U68/DATA1_10 , \U68/DATA1_11 ,
         \U63/DATA1_11 , \U58/DATA2_4 , \U58/DATA2_5 , \U58/DATA2_6 ,
         \U58/DATA2_7 , \U58/DATA2_8 , \U58/DATA2_9 , \U58/DATA1_4 ,
         \U58/DATA1_5 , \U58/DATA1_6 , \U58/DATA1_7 , \U58/DATA1_8 ,
         \U58/DATA1_9 , \U58/DATA1_10 , \U58/DATA1_11 , \U55/DATA2_11 ,
         \U55/DATA1_11 , \U50/DATA1_4 , \U50/DATA1_5 , \U50/DATA1_6 ,
         \U50/DATA1_7 , \U50/DATA1_8 , \U50/DATA1_9 , \U50/DATA1_10 ,
         \U50/DATA1_11 , \U45/DATA1_5 , \U45/DATA1_6 , \U45/DATA1_7 ,
         \U45/DATA1_8 , \U45/DATA1_9 , \U45/DATA1_10 , \U45/DATA1_11 ,
         \U40/DATA1_1 , \U40/DATA1_2 , \U40/DATA1_3 , \U40/DATA1_4 ,
         \U40/DATA1_5 , \U40/DATA1_6 , \U40/DATA1_7 , \U40/DATA1_8 ,
         \U40/DATA1_9 , \U40/DATA1_10 , \U40/DATA1_11 , \U35/DATA1_4 ,
         \U35/DATA1_5 , \U35/DATA1_6 , \U35/DATA1_7 , \U35/DATA1_8 ,
         \U35/DATA1_9 , \U35/DATA1_10 , \U35/DATA1_11 , \U30/DATA1_9 ,
         \U30/DATA1_10 , \U30/DATA1_11 , \U25/DATA1_1 , \U25/DATA1_2 ,
         \U25/DATA1_3 , \U25/DATA1_4 , \U25/DATA1_5 , \U25/DATA1_6 ,
         \U25/DATA1_7 , \U25/DATA1_8 , \U25/DATA1_9 , \U25/DATA1_10 ,
         \U25/DATA1_11 , \U20/DATA1_6 , \U20/DATA1_7 , \U20/DATA1_8 ,
         \U20/DATA1_9 , \U20/DATA1_10 , \U20/DATA1_11 , \U15/DATA1_11 ,
         \U10/DATA1_9 , \U10/DATA1_10 , \U10/DATA1_11 , \U5/DATA2_9 ,
         \U5/DATA1_9 , \U5/DATA1_10 , \U5/DATA1_11 , \U4/Z_9 , \U4/Z_10 ,
         \U4/Z_11 , \U4/Z_12 , \U4/Z_13 , \U4/Z_14 , \U4/Z_15 , \U4/Z_16 ,
         \U4/Z_17 , \U4/Z_18 , \U4/Z_19 , \U4/Z_20 , \U4/Z_21 , \U4/Z_22 ,
         \U4/Z_23 , \U4/Z_24 , \U4/Z_25 , \U4/Z_26 , \U4/Z_27 , \U4/Z_28 ,
         \U4/Z_29 , \U4/Z_30 , \U4/Z_31 , \U4/Z_32 , \U4/Z_33 , \U4/Z_34 ,
         \U4/Z_35 , \U4/Z_36 , \U4/Z_37 , \U4/Z_38 , \U4/Z_39 , \U4/Z_40 ,
         \U4/Z_41 , \U4/Z_42 , \U4/Z_43 , \U4/Z_44 , \U4/Z_45 , \U4/Z_46 ,
         \U4/Z_47 , \U4/Z_48 , \U4/Z_49 , \U4/Z_50 , \U4/Z_51 , \U4/Z_52 ,
         \U4/Z_53 , \U4/Z_54 , \fadd_0_0_0_0_0/syncressign_d1 ,
         \fadd_0_0_0_0_0/syncsigny_d2 , \fadd_0_0_0_0_0/syncsigny_d1 ,
         \fadd_0_0_0_0_0/synceffsub_d1 , \fadd_0_0_0_0_0/zerofromclose_d1 ,
         \fadd_0_0_0_0_0/zerofromclose , \fadd_0_0_0_0_0/round ,
         \fadd_0_0_0_0_0/expoperationsel[0] , \fadd_0_0_0_0_0/cinaddfar ,
         \fadd_0_0_0_0_0/ressign , \fadd_0_0_0_0_0/selectclosepath_d1 ,
         \fadd_0_0_0_0_0/effsub_d1 , \fadd_0_0_0_0_0/newy_9 ,
         \fadd_0_0_0_0_0/newy_10 , \fadd_0_0_0_0_0/newy_11 ,
         \fadd_0_0_0_0_1/syncressign_d1 , \fadd_0_0_0_0_1/syncsigny_d1 ,
         \fadd_0_0_0_0_1/synceffsub_d1 , \fadd_0_0_0_0_1/zerofromclose_d1 ,
         \fadd_0_0_0_0_1/zerofromclose , \fadd_0_0_0_0_1/round ,
         \fadd_0_0_0_0_1/expoperationsel[0] , \fadd_0_0_0_0_1/cinaddfar ,
         \fadd_0_0_0_0_1/ressign , \fadd_0_0_0_0_1/selectclosepath_d1 ,
         \fadd_0_0_0_0_1/effsub_d1 , \fadd_0_0_0_0_1/newy_9 ,
         \fadd_0_0_0_0_1/newy_10 , \fadd_0_0_0_0_1/newy_11 ,
         \fadd_0_0_0_0_2/syncressign_d1 , \fadd_0_0_0_0_2/syncsigny_d2 ,
         \fadd_0_0_0_0_2/syncsigny_d1 , \fadd_0_0_0_0_2/synceffsub_d1 ,
         \fadd_0_0_0_0_2/zerofromclose_d1 , \fadd_0_0_0_0_2/zerofromclose ,
         \fadd_0_0_0_0_2/round , \fadd_0_0_0_0_2/expoperationsel[0] ,
         \fadd_0_0_0_0_2/cinaddfar , \fadd_0_0_0_0_2/ressign ,
         \fadd_0_0_0_0_2/selectclosepath_d1 , \fadd_0_0_0_0_2/effsub_d1 ,
         \fadd_0_0_0_0_2/newy_9 , \fadd_0_0_0_0_2/newy_10 ,
         \fadd_0_0_0_0_2/newy_11 , \fadd_0_0_0_0_3/syncressign_d1 ,
         \fadd_0_0_0_0_3/syncsigny_d1 , \fadd_0_0_0_0_3/synceffsub_d1 ,
         \fadd_0_0_0_0_3/zerofromclose_d1 , \fadd_0_0_0_0_3/zerofromclose ,
         \fadd_0_0_0_0_3/round , \fadd_0_0_0_0_3/expoperationsel[0] ,
         \fadd_0_0_0_0_3/cinaddfar , \fadd_0_0_0_0_3/ressign ,
         \fadd_0_0_0_0_3/selectclosepath_d1 , \fadd_0_0_0_0_3/effsub_d1 ,
         \fadd_0_0_0_0_3/newy_9 , \fadd_0_0_0_0_3/newy_10 ,
         \fadd_0_0_0_0_3/newy_11 , \fadd_0_0_0_0_4/syncressign_d1 ,
         \fadd_0_0_0_0_4/syncsigny_d1 , \fadd_0_0_0_0_4/synceffsub_d1 ,
         \fadd_0_0_0_0_4/zerofromclose_d1 , \fadd_0_0_0_0_4/zerofromclose ,
         \fadd_0_0_0_0_4/round , \fadd_0_0_0_0_4/expoperationsel[0] ,
         \fadd_0_0_0_0_4/cinaddfar , \fadd_0_0_0_0_4/ressign ,
         \fadd_0_0_0_0_4/selectclosepath_d1 , \fadd_0_0_0_0_4/effsub_d1 ,
         \fadd_0_0_0_0_4/newy_9 , \fadd_0_0_0_0_4/newy_10 ,
         \fadd_0_0_0_0_4/newy_11 , \fadd_0_0_0_0_5/syncressign_d1 ,
         \fadd_0_0_0_0_5/syncsigny_d2 , \fadd_0_0_0_0_5/syncsigny_d1 ,
         \fadd_0_0_0_0_5/synceffsub_d1 , \fadd_0_0_0_0_5/zerofromclose_d1 ,
         \fadd_0_0_0_0_5/zerofromclose , \fadd_0_0_0_0_5/round ,
         \fadd_0_0_0_0_5/expoperationsel[0] , \fadd_0_0_0_0_5/cinaddfar ,
         \fadd_0_0_0_0_5/ressign , \fadd_0_0_0_0_5/selectclosepath_d1 ,
         \fadd_0_0_0_0_5/effsub_d1 , \fadd_0_0_0_0_5/newy_9 ,
         \fadd_0_0_0_0_5/newy_10 , \fadd_0_0_0_0_5/newy_11 ,
         \fadd_0_0_0_0_6/syncressign_d1 , \fadd_0_0_0_0_6/syncsigny_d2 ,
         \fadd_0_0_0_0_6/syncsigny_d1 , \fadd_0_0_0_0_6/synceffsub_d1 ,
         \fadd_0_0_0_0_6/zerofromclose_d1 , \fadd_0_0_0_0_6/zerofromclose ,
         \fadd_0_0_0_0_6/round , \fadd_0_0_0_0_6/expoperationsel[0] ,
         \fadd_0_0_0_0_6/cinaddfar , \fadd_0_0_0_0_6/ressign ,
         \fadd_0_0_0_0_6/selectclosepath_d1 , \fadd_0_0_0_0_6/effsub_d1 ,
         \fadd_0_0_0_0_6/newy_9 , \fadd_0_0_0_0_6/newy_10 ,
         \fadd_0_0_0_0_6/newy_11 , \fadd_0_0_0_0_7/syncressign_d1 ,
         \fadd_0_0_0_0_7/syncsigny_d2 , \fadd_0_0_0_0_7/syncsigny_d1 ,
         \fadd_0_0_0_0_7/synceffsub_d1 , \fadd_0_0_0_0_7/zerofromclose_d1 ,
         \fadd_0_0_0_0_7/zerofromclose , \fadd_0_0_0_0_7/round ,
         \fadd_0_0_0_0_7/expoperationsel[0] , \fadd_0_0_0_0_7/cinaddfar ,
         \fadd_0_0_0_0_7/ressign , \fadd_0_0_0_0_7/selectclosepath_d1 ,
         \fadd_0_0_0_0_7/effsub_d1 , \fadd_0_0_0_0_7/newy_9 ,
         \fadd_0_0_0_0_7/newy_10 , \fadd_0_0_0_0_7/newy_11 ,
         \fadd_0_0_0_0_8/syncressign_d1 , \fadd_0_0_0_0_8/syncsigny_d1 ,
         \fadd_0_0_0_0_8/synceffsub_d1 , \fadd_0_0_0_0_8/zerofromclose_d1 ,
         \fadd_0_0_0_0_8/zerofromclose , \fadd_0_0_0_0_8/round ,
         \fadd_0_0_0_0_8/expoperationsel[0] , \fadd_0_0_0_0_8/cinaddfar ,
         \fadd_0_0_0_0_8/ressign , \fadd_0_0_0_0_8/selectclosepath_d1 ,
         \fadd_0_0_0_0_8/effsub_d1 , \fadd_0_0_0_0_8/newy_9 ,
         \fadd_0_0_0_0_8/newy_10 , \fadd_0_0_0_0_8/newy_11 ,
         \fadd_0_0_0_0_9/syncressign_d1 , \fadd_0_0_0_0_9/syncsigny_d1 ,
         \fadd_0_0_0_0_9/synceffsub_d1 , \fadd_0_0_0_0_9/zerofromclose_d1 ,
         \fadd_0_0_0_0_9/zerofromclose , \fadd_0_0_0_0_9/round ,
         \fadd_0_0_0_0_9/expoperationsel[0] , \fadd_0_0_0_0_9/cinaddfar ,
         \fadd_0_0_0_0_9/ressign , \fadd_0_0_0_0_9/selectclosepath_d1 ,
         \fadd_0_0_0_0_9/effsub_d1 , \fadd_0_0_0_0_9/newy_9 ,
         \fadd_0_0_0_0_9/newy_10 , \fadd_0_0_0_0_9/newy_11 ,
         \fadd_0_0_0_0_10/sub_707/carry[5] ,
         \fadd_0_0_0_0_10/sub_707/carry[4] ,
         \fadd_0_0_0_0_10/sub_707/carry[3] ,
         \fadd_0_0_0_0_10/sub_707/carry[2] ,
         \fadd_0_0_0_0_10/sub_707/carry[1] ,
         \fadd_0_0_0_0_10/sub_710/carry[4] ,
         \fadd_0_0_0_0_10/sub_710/carry[3] ,
         \fadd_0_0_0_0_10/sub_710/carry[2] ,
         \fadd_0_0_0_0_10/sub_710/carry[1] , \fadd_0_0_0_0_10/sub_784/A[2] ,
         \fadd_0_0_0_0_10/sub_784/A[1] , \fadd_0_0_0_0_10/sub_784/DIFF[4] ,
         \fadd_0_0_0_0_10/sub_784/DIFF[3] , \fadd_0_0_0_0_10/sub_784/DIFF[2] ,
         \fadd_0_0_0_0_10/sub_784/DIFF[1] , \fadd_0_0_0_0_10/sub_784/DIFF[0] ,
         \fadd_0_0_0_0_10/sub_784/carry[4] ,
         \fadd_0_0_0_0_10/sub_784/carry[3] ,
         \fadd_0_0_0_0_10/sub_784/carry[2] ,
         \fadd_0_0_0_0_10/sub_784/carry[1] ,
         \fadd_0_0_0_0_10/add_859/carry[6] , \fadd_0_0_0_0_10/U4/DATA1_10 ,
         \fadd_0_0_0_0_10/U4/DATA1_9 , \fadd_0_0_0_0_10/U4/DATA1_7 ,
         \fadd_0_0_0_0_10/U4/DATA1_6 , \fadd_0_0_0_0_10/U4/DATA1_4 ,
         \fadd_0_0_0_0_10/U4/DATA2_10 , \fadd_0_0_0_0_10/U5/DATA1_4 ,
         \fadd_0_0_0_0_10/U5/DATA1_3 , \fadd_0_0_0_0_10/U5/DATA1_2 ,
         \fadd_0_0_0_0_10/U5/DATA1_1 , \fadd_0_0_0_0_10/U5/DATA1_0 ,
         \fadd_0_0_0_0_10/U5/DATA2_4 , \fadd_0_0_0_0_10/U5/DATA2_3 ,
         \fadd_0_0_0_0_10/U5/DATA2_2 , \fadd_0_0_0_0_10/U5/DATA2_1 ,
         \fadd_0_0_0_0_10/U5/DATA2_0 , \fadd_0_0_0_0_10/U11/DATA2_8 ,
         \fadd_0_0_0_0_10/U11/DATA2_7 , \fadd_0_0_0_0_10/U11/DATA2_6 ,
         \fadd_0_0_0_0_10/U11/DATA2_5 , \fadd_0_0_0_0_10/U11/DATA2_3 ,
         \fadd_0_0_0_0_10/U11/DATA2_2 , \fadd_0_0_0_0_10/U11/DATA2_1 ,
         \fadd_0_0_0_0_10/U11/DATA2_0 , \fadd_0_0_0_0_10/U12/DATA3_0 ,
         \fadd_0_0_0_0_10/U20/DATA1_0 , \fadd_0_0_0_0_10/U21/DATA2_3 ,
         \fadd_0_0_0_0_10/U21/DATA2_2 , \fadd_0_0_0_0_10/U22/DATA1_3 ,
         \fadd_0_0_0_0_10/U22/DATA1_2 , \fadd_0_0_0_0_10/U22/DATA1_1 ,
         \fadd_0_0_0_0_10/U22/DATA1_0 , \fadd_0_0_0_0_10/U23/Z_0 ,
         \fadd_0_0_0_0_10/U24/DATA1_5 , \fadd_0_0_0_0_10/U24/DATA1_4 ,
         \fadd_0_0_0_0_10/U24/DATA1_3 , \fadd_0_0_0_0_10/U24/DATA1_2 ,
         \fadd_0_0_0_0_10/U24/DATA1_1 , \fadd_0_0_0_0_10/U24/DATA2_5 ,
         \fadd_0_0_0_0_10/U24/DATA2_4 , \fadd_0_0_0_0_10/U24/DATA2_3 ,
         \fadd_0_0_0_0_10/U24/DATA2_2 , \fadd_0_0_0_0_10/U24/DATA2_1 ,
         \fadd_0_0_0_0_10/U24/Z_5 , \fadd_0_0_0_0_10/U24/Z_4 ,
         \fadd_0_0_0_0_10/U24/Z_3 , \fadd_0_0_0_0_10/U24/Z_2 ,
         \fadd_0_0_0_0_10/U24/Z_1 , \fadd_0_0_0_0_10/U25/Z_3 ,
         \fadd_0_0_0_0_10/U25/Z_2 , \fadd_0_0_0_0_10/U27/DATA1_0 ,
         \fadd_0_0_0_0_10/U27/Z_2 , \fadd_0_0_0_0_10/U27/Z_1 ,
         \fadd_0_0_0_0_10/U28/Z_6 , \fadd_0_0_0_0_10/U28/Z_5 ,
         \fadd_0_0_0_0_10/U28/Z_4 , \fadd_0_0_0_0_10/U29/Z_11 ,
         \fadd_0_0_0_0_10/U29/Z_10 , \fadd_0_0_0_0_10/U29/Z_8 ,
         \fadd_0_0_0_0_10/U29/Z_7 , \fadd_0_0_0_0_10/U29/Z_6 ,
         \fadd_0_0_0_0_10/U29/Z_5 , \fadd_0_0_0_0_10/U29/Z_4 ,
         \fadd_0_0_0_0_10/U29/Z_3 , \fadd_0_0_0_0_10/U29/Z_2 ,
         \fadd_0_0_0_0_10/U29/Z_1 , \fadd_0_0_0_0_10/U29/Z_0 ,
         \fadd_0_0_0_0_10/n305 , \fadd_0_0_0_0_10/n302 ,
         \fadd_0_0_0_0_10/n240 , \fadd_0_0_0_0_10/n239 ,
         \fadd_0_0_0_0_10/n238 , \fadd_0_0_0_0_10/n237 ,
         \fadd_0_0_0_0_10/n236 , \fadd_0_0_0_0_10/n235 ,
         \fadd_0_0_0_0_10/n234 , \fadd_0_0_0_0_10/n213 ,
         \fadd_0_0_0_0_10/n212 , \fadd_0_0_0_0_10/n211 ,
         \fadd_0_0_0_0_10/n210 , \fadd_0_0_0_0_10/n209 ,
         \fadd_0_0_0_0_10/n182 , \fadd_0_0_0_0_10/n169 ,
         \fadd_0_0_0_0_10/n168 , \fadd_0_0_0_0_10/n167 ,
         \fadd_0_0_0_0_10/n166 , \fadd_0_0_0_0_10/n165 ,
         \fadd_0_0_0_0_10/n164 , \fadd_0_0_0_0_10/n163 ,
         \fadd_0_0_0_0_10/n162 , \fadd_0_0_0_0_10/n161 ,
         \fadd_0_0_0_0_10/n160 , \fadd_0_0_0_0_10/n159 ,
         \fadd_0_0_0_0_10/n148 , \fadd_0_0_0_0_10/n147 ,
         \fadd_0_0_0_0_10/n146 , \fadd_0_0_0_0_10/n145 ,
         \fadd_0_0_0_0_10/n144 , \fadd_0_0_0_0_10/n143 ,
         \fadd_0_0_0_0_10/n142 ,
         \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_dualsubclose/sub_1_root_add_300/carry[6] ,
         \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_dualsubclose/sub_1_root_add_300/carry[5] ,
         \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_dualsubclose/sub_1_root_add_300/carry[4] ,
         \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_dualsubclose/sub_1_root_add_300/carry[3] ,
         \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_dualsubclose/sub_1_root_add_300/carry[2] ,
         \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_dualsubclose/sub_1_root_add_303/carry[5] ,
         \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_dualsubclose/sub_1_root_add_303/carry[4] ,
         \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_dualsubclose/sub_1_root_add_303/carry[3] ,
         \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_dualsubclose/sub_1_root_add_303/carry[2] ,
         \fadd_0_0_0_0_0/norm/level1_d1[4] ,
         \fadd_0_0_0_0_1/norm/level1_d1[4] ,
         \fadd_0_0_0_0_2/norm/level1_d1[4] ,
         \fadd_0_0_0_0_3/norm/level1_d1[4] ,
         \fadd_0_0_0_0_4/norm/level1_d1[4] ,
         \fadd_0_0_0_0_5/norm/level1_d1[4] ,
         \fadd_0_0_0_0_6/norm/level1_d1[4] ,
         \fadd_0_0_0_0_7/norm/level1_d1[4] ,
         \fadd_0_0_0_0_8/norm/level1_d1[4] ,
         \fadd_0_0_0_0_9/norm/level1_d1[4] , \fadd_0_0_0_0_10/norm/U4/DATA2_5 ,
         \fadd_0_0_0_0_10/norm/U5/Z_5 , \fadd_0_0_0_0_10/norm/U5/Z_4 ,
         \fadd_0_0_0_0_10/norm/U5/Z_3 , \fadd_0_0_0_0_10/norm/U5/Z_2 ,
         \fadd_0_0_0_0_10/norm/U5/Z_1 , \fadd_0_0_0_0_10/norm/U5/Z_0 ,
         \fadd_0_0_0_0_0/rightshiftercomponent/n389_o ,
         \fadd_0_0_0_0_0/rightshiftercomponent/level1_d2[0] ,
         \fadd_0_0_0_0_0/rightshiftercomponent/level1_d1[0] ,
         \fadd_0_0_0_0_0/rightshiftercomponent/level2[1] ,
         \fadd_0_0_0_0_0/rightshiftercomponent/ps_d2[0] ,
         \fadd_0_0_0_0_1/rightshiftercomponent/n389_o ,
         \fadd_0_0_0_0_1/rightshiftercomponent/level1_d2[0] ,
         \fadd_0_0_0_0_1/rightshiftercomponent/level1_d1[0] ,
         \fadd_0_0_0_0_1/rightshiftercomponent/level2[1] ,
         \fadd_0_0_0_0_1/rightshiftercomponent/ps_d2[0] ,
         \fadd_0_0_0_0_2/rightshiftercomponent/n389_o ,
         \fadd_0_0_0_0_2/rightshiftercomponent/level1_d2[0] ,
         \fadd_0_0_0_0_2/rightshiftercomponent/level1_d1[0] ,
         \fadd_0_0_0_0_2/rightshiftercomponent/level2[1] ,
         \fadd_0_0_0_0_2/rightshiftercomponent/ps_d2[0] ,
         \fadd_0_0_0_0_3/rightshiftercomponent/n389_o ,
         \fadd_0_0_0_0_3/rightshiftercomponent/level1_d2[0] ,
         \fadd_0_0_0_0_3/rightshiftercomponent/level1_d1[0] ,
         \fadd_0_0_0_0_3/rightshiftercomponent/level2[1] ,
         \fadd_0_0_0_0_3/rightshiftercomponent/ps_d2[0] ,
         \fadd_0_0_0_0_4/rightshiftercomponent/n389_o ,
         \fadd_0_0_0_0_4/rightshiftercomponent/level1_d2[0] ,
         \fadd_0_0_0_0_4/rightshiftercomponent/level1_d1[0] ,
         \fadd_0_0_0_0_4/rightshiftercomponent/level2[1] ,
         \fadd_0_0_0_0_4/rightshiftercomponent/ps_d2[0] ,
         \fadd_0_0_0_0_5/rightshiftercomponent/n389_o ,
         \fadd_0_0_0_0_5/rightshiftercomponent/level1_d2[0] ,
         \fadd_0_0_0_0_5/rightshiftercomponent/level1_d1[0] ,
         \fadd_0_0_0_0_5/rightshiftercomponent/level2[1] ,
         \fadd_0_0_0_0_5/rightshiftercomponent/ps_d2[0] ,
         \fadd_0_0_0_0_6/rightshiftercomponent/n389_o ,
         \fadd_0_0_0_0_6/rightshiftercomponent/level1_d2[0] ,
         \fadd_0_0_0_0_6/rightshiftercomponent/level1_d1[0] ,
         \fadd_0_0_0_0_6/rightshiftercomponent/level2[1] ,
         \fadd_0_0_0_0_6/rightshiftercomponent/ps_d2[0] ,
         \fadd_0_0_0_0_7/rightshiftercomponent/n389_o ,
         \fadd_0_0_0_0_7/rightshiftercomponent/level1_d2[0] ,
         \fadd_0_0_0_0_7/rightshiftercomponent/level1_d1[0] ,
         \fadd_0_0_0_0_7/rightshiftercomponent/level2[1] ,
         \fadd_0_0_0_0_7/rightshiftercomponent/ps_d2[0] ,
         \fadd_0_0_0_0_8/rightshiftercomponent/n389_o ,
         \fadd_0_0_0_0_8/rightshiftercomponent/level1_d2[0] ,
         \fadd_0_0_0_0_8/rightshiftercomponent/level1_d1[0] ,
         \fadd_0_0_0_0_8/rightshiftercomponent/level2[1] ,
         \fadd_0_0_0_0_8/rightshiftercomponent/ps_d2[0] ,
         \fadd_0_0_0_0_9/rightshiftercomponent/n389_o ,
         \fadd_0_0_0_0_9/rightshiftercomponent/level1_d2[0] ,
         \fadd_0_0_0_0_9/rightshiftercomponent/level1_d1[0] ,
         \fadd_0_0_0_0_9/rightshiftercomponent/level2[1] ,
         \fadd_0_0_0_0_9/rightshiftercomponent/ps_d2[0] ,
         \fadd_0_0_0_0_10/rightshiftercomponent/U5/Z_0 ,
         \fadd_0_0_0_0_10/rightshiftercomponent/U6/Z_0 ,
         \fadd_0_0_0_0_10/rightshiftercomponent/n44 ,
         \fadd_0_0_0_0_10/rightshiftercomponent/n43 ,
         \fadd_0_0_0_0_10/rightshiftercomponent/n42 ,
         \fadd_0_0_0_0_10/rightshiftercomponent/n41 ,
         \fadd_0_0_0_0_10/rightshiftercomponent/n17 ,
         \fadd_0_0_0_0_10/rightshiftercomponent/n16 ,
         \fadd_0_0_0_0_10/rightshiftercomponent/n11 ,
         \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/A[5] ,
         \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/A[4] ,
         \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/A[3] ,
         \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/A[2] ,
         \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/B[7] ,
         \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/B[6] ,
         \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/B[5] ,
         \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/B[4] ,
         \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/B[3] ,
         \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/B[2] ,
         \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/B[1] ,
         \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/B[0] ,
         \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/CI ,
         \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/SUM[7] ,
         \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/carry[7] ,
         \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/carry[6] ,
         \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/carry[5] ,
         \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/carry[4] ,
         \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/carry[3] ,
         \fmul_0_0_0_0_0/round , \fmul_0_0_0_0_0/sign , \fmul_0_0_0_0_1/round ,
         \fmul_0_0_0_0_1/sign , \fmul_0_0_0_0_2/round , \fmul_0_0_0_0_2/sign ,
         \fmul_0_0_0_0_3/round , \fmul_0_0_0_0_3/sign , \fmul_0_0_0_0_4/round ,
         \fmul_0_0_0_0_4/sign , \fmul_0_0_0_0_5/round , \fmul_0_0_0_0_5/sign ,
         \fmul_0_0_0_0_6/round , \fmul_0_0_0_0_6/sign , \fmul_0_0_0_0_7/round ,
         \fmul_0_0_0_0_7/sign , \fmul_0_0_0_0_8/expsigpostround[10] ,
         \fmul_0_0_0_0_8/round , \fmul_0_0_0_0_8/sign , \fmul_0_0_0_0_9/round ,
         \fmul_0_0_0_0_9/sign , \fmul_0_0_0_0_10/add_2_root_add_321/A[4] ,
         \fmul_0_0_0_0_10/add_2_root_add_321/A[3] ,
         \fmul_0_0_0_0_10/add_2_root_add_321/A[2] ,
         \fmul_0_0_0_0_10/add_2_root_add_321/A[1] ,
         \fmul_0_0_0_0_10/add_2_root_add_321/A[0] ,
         \fmul_0_0_0_0_10/add_2_root_add_321/B[4] ,
         \fmul_0_0_0_0_10/add_2_root_add_321/B[3] ,
         \fmul_0_0_0_0_10/add_2_root_add_321/B[2] ,
         \fmul_0_0_0_0_10/add_2_root_add_321/B[1] ,
         \fmul_0_0_0_0_10/add_2_root_add_321/B[0] ,
         \fmul_0_0_0_0_10/add_2_root_add_321/carry[5] ,
         \fmul_0_0_0_0_10/add_2_root_add_321/carry[4] ,
         \fmul_0_0_0_0_10/add_2_root_add_321/carry[3] ,
         \fmul_0_0_0_0_10/add_2_root_add_321/carry[2] ,
         \fmul_0_0_0_0_10/add_2_root_add_321/carry[1] ,
         \fmul_0_0_0_0_10/sub_1_root_add_321/A[4] ,
         \fmul_0_0_0_0_10/sub_1_root_add_321/A[3] ,
         \fmul_0_0_0_0_10/sub_1_root_add_321/A[2] ,
         \fmul_0_0_0_0_10/sub_1_root_add_321/A[1] ,
         \fmul_0_0_0_0_10/sub_1_root_add_321/A[0] ,
         \fmul_0_0_0_0_10/sub_1_root_add_321/DIFF[5] ,
         \fmul_0_0_0_0_10/sub_1_root_add_321/DIFF[4] ,
         \fmul_0_0_0_0_10/sub_1_root_add_321/DIFF[3] ,
         \fmul_0_0_0_0_10/sub_1_root_add_321/DIFF[2] ,
         \fmul_0_0_0_0_10/sub_1_root_add_321/DIFF[1] ,
         \fmul_0_0_0_0_10/sub_1_root_add_321/carry[5] ,
         \fmul_0_0_0_0_10/U8/Z_8 , \fmul_0_0_0_0_10/U8/Z_7 ,
         \fmul_0_0_0_0_10/U8/Z_6 , \fmul_0_0_0_0_10/U8/Z_5 ,
         \fmul_0_0_0_0_10/U9/Z_1 , \fmul_0_0_0_0_10/U9/Z_0 ,
         \fmul_0_0_0_0_10/n137 , \fmul_0_0_0_0_10/n98 ,
         \fmul_0_0_0_0_0/roundingadder/n151_o[0] ,
         \fmul_0_0_0_0_1/roundingadder/n151_o[0] ,
         \fmul_0_0_0_0_2/roundingadder/n151_o[0] ,
         \fmul_0_0_0_0_3/roundingadder/n151_o[0] ,
         \fmul_0_0_0_0_4/roundingadder/n151_o[0] ,
         \fmul_0_0_0_0_5/roundingadder/n151_o[0] ,
         \fmul_0_0_0_0_6/roundingadder/n151_o[0] ,
         \fmul_0_0_0_0_7/roundingadder/n151_o[0] ,
         \fmul_0_0_0_0_8/roundingadder/n151_o[0] ,
         \fmul_0_0_0_0_9/roundingadder/n151_o[0] ,
         \fmul_0_0_0_0_10/roundingadder/add_1_root_add_57/A[9] ,
         \fmul_0_0_0_0_10/roundingadder/add_1_root_add_57/A[8] ,
         \fmul_0_0_0_0_10/roundingadder/add_1_root_add_57/A[7] ,
         \fmul_0_0_0_0_10/roundingadder/add_1_root_add_57/A[6] ,
         \fmul_0_0_0_0_10/roundingadder/add_1_root_add_57/A[5] ,
         \fmul_0_0_0_0_10/roundingadder/add_1_root_add_57/A[4] ,
         \fmul_0_0_0_0_10/roundingadder/add_1_root_add_57/A[3] ,
         \fmul_0_0_0_0_10/roundingadder/add_1_root_add_57/A[2] ,
         \fmul_0_0_0_0_10/roundingadder/add_1_root_add_57/A[1] ,
         \fmul_0_0_0_0_10/roundingadder/add_1_root_add_57/A[0] ,
         \fmul_0_0_0_0_10/roundingadder/add_1_root_add_57/CI ,
         \fmul_0_0_0_0_10/roundingadder/add_1_root_add_57/SUM[10] ,
         \fmul_0_0_0_0_10/roundingadder/add_1_root_add_57/SUM[9] , n8208,
         n8216, n8219, n8222, n8225, n8228, n8231, n8234, n8237, n8240, n8245,
         n8247, n8250, n8254, n8258, n8262, n8266, n8270, n8274, n8278, n8282,
         n8285, n8289, n8292, n8295, n8298, n8301, n8304, n8307, n8310, n8313,
         n8316, n8319, n8322, n8325, n8328, n8331, n8336, n8340, n8344, n8348,
         n8352, n8356, n8360, n8364, n8368, n8372, n8376, n8380, n8383, n8386,
         n8389, n8392, n8395, n8398, n8401, n8404, n8407, n8416, n8419, n8422,
         n8425, n8428, n8431, n8434, n8437, n8440, n8443, n8446, n8449, n8452,
         n8455, n8458, n8461, n8464, n8467, n8470, n8473, n8476, n8479, n8482,
         n8485, n8488, n8491, n8494, n8497, n8500, n8503, n8506, n8509, n8512,
         n8515, n8518, n8521, n8523, n8527, n8530, n8533, n8536, n8539, n8542,
         n8545, n8548, n8551, n8557, n8560, n8563, n8566, n8569, n8572, n8575,
         n8578, n8581, n8584, n8587, n8590, n8593, n8596, n8599, n8602, n8605,
         n8608, n8611, n8614, n8617, n8620, n8623, n8626, n8629, n8632, n8633,
         n8636, n8637, n8640, n8641, n8644, n8645, n8648, n8649, n8652, n8653,
         n8656, n8657, n8660, n8661, n8664, n8665, n8668, n8669, n8671, n8672,
         n8673, n8674, n8678, n8679, n8680, n8681, n8682, n8683, n8685, n8686,
         n8687, n8689, n8690, n8691, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8713, n8714, n8715, n8716, n8717, n8723, n8724, n8725,
         n8726, n8730, n8731, n8732, n8734, n8735, n8738, n8739, n8741, n8742,
         n8744, n8745, n8747, n8748, n8750, n8751, n8753, n8754, n8756, n8757,
         n8759, n8760, n8763, n8764, n8766, n8768, n8770, n8771, n8774, n8776,
         n8777, n8778, n8780, n8781, n8782, n8784, n8787, n8789, n8790, n8791,
         n8793, n8794, n8796, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8808, n8809, n8810, n8811, n8812, n8814, n8815, n8817, n8818,
         n8819, n8822, n8823, n8824, n8826, n8827, n8828, n8830, n8831, n8833,
         n8834, n8836, n8837, n8838, n8839, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8849, n8850, n8852, n8853, n8854, n8855, n8856, n8860,
         n8861, n8862, n8863, n8866, n8867, n8869, n8870, n8871, n8873, n8874,
         n8875, n8877, n8878, n8879, n8881, n8882, n8883, n8884, n8886, n8887,
         n8893, n8894, n8906, n8910, n8912, n8915, n8916, n8917, n8929, n8935,
         n8936, n8947, n8949, n8953, n8955, n8958, n8960, n8961, n8964, n8965,
         n8967, n8968, n8970, n8972, n8974, n8976, n8978, n8980, n8982, n8984,
         n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9007, n9008, n9009, n9010, n9011,
         n9012, n9016, n9017, n9021, n9022, n9026, n9027, n9031, n9032, n9036,
         n9037, n9041, n9042, n9046, n9047, n9051, n9052, n9055, n9057, n9058,
         n9060, n9062, n9065, n9066, n9068, n9070, n9071, n9074, n9075, n9076,
         n9078, n9080, n9082, n9084, n9086, n9088, n9090, n9092, n9094, n9096,
         n9097, n9099, n9100, n9102, n9106, n9107, n9108, n9110, n9112, n9114,
         n9116, n9118, n9120, n9122, n9124, n9126, n9128, n9129, n9130, n9132,
         n9134, n9136, n9139, n9141, n9142, n9144, n9145, n9147, n9148, n9150,
         n9152, n9154, n9156, n9158, n9160, n9162, n9164, n9166, n9167, n9168,
         n9171, n9174, n9175, n9177, n9178, n9179, n9181, n9183, n9185, n9187,
         n9189, n9191, n9193, n9195, n9198, n9202, n9204, n9207, n9208, n9210,
         n9221, n9227, n9228, n9240, n9244, n9246, n9249, n9250, n9252, n9263,
         n9269, n9270, n9281, n9285, n9286, n9288, n9290, n9291, n9293, n9294,
         n9296, n9297, n9299, n9301, n9303, n9305, n9307, n9309, n9311, n9313,
         n9315, n9316, n9319, n9322, n9323, n9325, n9326, n9327, n9329, n9331,
         n9333, n9335, n9337, n9339, n9341, n9343, n9346, n9350, n9352, n9355,
         n9356, n9357, n9369, n9375, n9376, n9388, n9392, n9394, n9397, n9398,
         n9399, n9410, n9412, n9418, n9419, n9430, n9431, n9436, n9439, n9440,
         n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9450, n9451,
         n9452, n9453, n9454, n9455, n9457, n9458, n9459, n9460, n9461, n9462,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9501, n9502, n9503, n9504,
         n9505, n9506, n9508, n9509, n9510, n9511, n9512, n9513, n9515, n9516,
         n9517, n9518, n9519, n9520, n9522, n9523, n9524, n9525, n9526, n9527,
         n9529, n9531, n9533, n9534, n9535, n9536, n9537, n9538, n9540, n9542,
         n9544, n9546, n9547, n9548, n9549, n9550, n9551, n9553, n9554, n9555,
         n9556, n9557, n9558, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
         n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
         n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
         n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
         n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606,
         n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
         n9617, n9618, n9619, n9624, n9625, n9626, n9627, n9628, n9629, n9631,
         n9632, n9633, n9634, n9635, n9636, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9702, n9703, n9704, n9705, n9706,
         n9707, n9709, n9710, n9711, n9712, n9713, n9714, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9780, n9781, n9782,
         n9783, n9784, n9785, n9787, n9788, n9789, n9790, n9791, n9792, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9858,
         n9859, n9860, n9861, n9862, n9863, n9865, n9866, n9867, n9868, n9869,
         n9870, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9936, n9937, n9938, n9939, n9940, n9941, n9943, n9944, n9945,
         n9946, n9947, n9948, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10014, n10015, n10016, n10017,
         n10018, n10019, n10021, n10022, n10023, n10024, n10025, n10026,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10092, n10093, n10094, n10095,
         n10096, n10097, n10099, n10100, n10101, n10102, n10103, n10104,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10170, n10171, n10172, n10173,
         n10174, n10175, n10177, n10178, n10179, n10180, n10181, n10182,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10248, n10249, n10250, n10251,
         n10252, n10253, n10255, n10256, n10257, n10258, n10259, n10260,
         n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
         n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
         n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
         n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
         n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301,
         n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309,
         n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317,
         n10318, n10319, n10320, n10321, n10323, n10324, n10325, n10326,
         n10327, n10328, n10330, n10331, n10332, n10333, n10334, n10335,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10399, n10400, n10402,
         n10404, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10446, n10447, n10448, n10449, n10450, n10451, n10452,
         n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10462,
         n10463, n10464, n10465, n10466, n10467, n10468, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10502, n10503, n10505, n10506,
         n10507, n10509, n10510, n10511, n10512, n10513, n10514, n10515,
         n10516, n10517, n10518, n10519, n10521, n10522, n10523, n10524,
         n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532,
         n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540,
         n10541, n10542, n10544, n10545, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10586, n10587,
         n10588, n10592, n10593, n10594, n10596, n10597, n10599, n10601,
         n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
         n10611, n10612, n10613, n10614, n10616, n10617, n10620, n10625,
         n10626, n10627, n10630, n10632, n10633, n10634, n10635, n10636,
         n10637, n10638, n10640, n10642, n10643, n10644, n10645, n10646,
         n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654,
         n10655, n10656, n10657, n10658, n10663, n10664, n10667, n10668,
         n10669, n10673, n10674, n10675, n10677, n10678, n10680, n10682,
         n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691,
         n10692, n10693, n10694, n10695, n10697, n10698, n10701, n10706,
         n10707, n10710, n10713, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10723, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10746, n10747, n10750, n10751,
         n10752, n10756, n10757, n10758, n10760, n10761, n10763, n10765,
         n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774,
         n10775, n10776, n10777, n10778, n10780, n10781, n10784, n10789,
         n10790, n10791, n10794, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10804, n10806, n10807, n10808, n10809, n10810,
         n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818,
         n10819, n10820, n10821, n10822, n10827, n10828, n10831, n10832,
         n10833, n10837, n10838, n10839, n10841, n10842, n10844, n10846,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10861, n10862, n10865, n10870,
         n10871, n10872, n10875, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10885, n10887, n10888, n10889, n10890, n10891,
         n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899,
         n10900, n10901, n10902, n10903, n10908, n10909, n10912, n10913,
         n10914, n10918, n10919, n10920, n10922, n10923, n10925, n10927,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10942, n10943, n10946, n10951,
         n10952, n10953, n10956, n10958, n10959, n10960, n10961, n10962,
         n10963, n10964, n10966, n10968, n10969, n10970, n10971, n10972,
         n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980,
         n10981, n10982, n10983, n10984, n10989, n10990, n10993, n10994,
         n10995, n10999, n11000, n11001, n11003, n11004, n11006, n11008,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11023, n11024, n11027, n11032,
         n11033, n11034, n11037, n11039, n11040, n11041, n11042, n11043,
         n11044, n11045, n11047, n11049, n11050, n11051, n11052, n11053,
         n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061,
         n11062, n11063, n11064, n11065, n11070, n11071, n11074, n11075,
         n11076, n11080, n11081, n11082, n11084, n11085, n11087, n11089,
         n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,
         n11099, n11100, n11101, n11102, n11104, n11105, n11108, n11113,
         n11114, n11115, n11118, n11120, n11121, n11122, n11123, n11124,
         n11125, n11126, n11128, n11130, n11131, n11132, n11133, n11134,
         n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142,
         n11143, n11144, n11145, n11146, n11151, n11152, n11155, n11156,
         n11157, n11161, n11162, n11163, n11165, n11166, n11168, n11170,
         n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179,
         n11180, n11181, n11182, n11183, n11185, n11186, n11189, n11194,
         n11195, n11196, n11199, n11201, n11202, n11203, n11204, n11205,
         n11206, n11207, n11209, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11232, n11233, n11234, n11235,
         n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
         n11245, n11246, n11247, n11249, n11250, n11251, n11252, n11253,
         n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11262,
         n11263, n11264, n11266, n11267, n11268, n11271, n11272, n11273,
         n11275, n11276, n11277, n11279, n11280, n11281, n11282, n11283,
         n11284, n11285, n11286, n11287, n11288, n11291, n11292, n11293,
         n11297, n11298, n11299, n11301, n11302, n11304, n11306, n11308,
         n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316,
         n11317, n11318, n11319, n11321, n11322, n11325, n11330, n11331,
         n11332, n11335, n11337, n11338, n11339, n11340, n11341, n11342,
         n11343, n11345, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11368, n11369, n11372, n11373, n11374,
         n11378, n11379, n11380, n11382, n11383, n11385, n11387, n11389,
         n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397,
         n11398, n11399, n11400, n11402, n11403, n11406, n11411, n11412,
         n11415, n11418, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11428, n11430, n11431, n11432, n11433, n11434, n11435,
         n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
         n11444, n11445, n11446, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11470, n11471, n11472,
         n11476, n11477, n11478, n11479, n11481, n11483, n11484, n11485,
         n11489, n11490, n11491, n11492, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11505, n11506,
         n11507, n11511, n11512, n11513, n11514, n11516, n11518, n11519,
         n11520, n11524, n11525, n11526, n11527, n11529, n11531, n11532,
         n11533, n11537, n11538, n11539, n11540, n11542, n11544, n11545,
         n11546, n11550, n11551, n11552, n11553, n11555, n11557, n11558,
         n11559, n11563, n11564, n11565, n11566, n11568, n11570, n11571,
         n11572, n11576, n11577, n11578, n11579, n11581, n11583, n11584,
         n11585, n11589, n11590, n11591, n11592, n11594, n11596, n11597,
         n11598, n11602, n11603, n11604, n11605, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11665, n11666, n11667, n11668, n11669, n11670,
         n11676, n11677, n11678, n11679, n11680, n11686, n11687, n11688,
         n11689, n11690, n11691, n11697, n11698, n11699, n11700, n11701,
         n11707, n11708, n11709, n11710, n11711, n11712, n11718, n11719,
         n11720, n11721, n11722, n11728, n11729, n11730, n11731, n11732,
         n11733, n11739, n11740, n11741, n11742, n11743, n11749, n11750,
         n11751, n11752, n11753, n11754, n11760, n11761, n11762, n11763,
         n11764, n11770, n11771, n11772, n11773, n11774, n11775, n11781,
         n11782, n11783, n11784, n11785, n11791, n11792, n11793, n11794,
         n11795, n11796, n11802, n11803, n11804, n11805, n11806, n11812,
         n11813, n11814, n11815, n11816, n11817, n11823, n11824, n11825,
         n11826, n11827, n11833, n11834, n11835, n11836, n11837, n11838,
         n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851,
         n11852, n11853, n11854, n11856, n11857, n11858, n11859, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11877, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11939, n11941, n11943, n11945, n11947, n11949, n11951, n11952,
         n11953, n11954, n11956, n11958, n11959, n11960, n11961, n11963,
         n11964, n11965, n11967, n11968, n11969, n11971, n11972, n11973,
         n11975, n11976, n11977, n11979, n11980, n11981, n11983, n11984,
         n11985, n11987, n11988, n11989, n11991, n11992, n11993, n11995,
         n11996, n11997, n11999, n12000, n12001, n12002, n12004, n12005,
         n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013,
         n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12024,
         n12028, n12032, n12036, n12037, n12041, n12042, n12055, n12056,
         n12057, n12061, n12062, n12063, n12065, n12066, n12067, n12068,
         n12069, n12070, n12071, n12072, n12073, n12094, n12095, n12097,
         n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12107,
         n12109, n12111, n12114, n12117, n12120, n12123, n12126, n12129,
         n12132, n12135, n12138, n12140, n12142, n12143, n12146, n12147,
         n12148, n12169, n12174, n12175, n12176, n12177, n12178, n12179,
         n12181, n12182, n12203, n12207, n12208, n12209, n12211, n12212,
         n12231, n12237, n12238, n12239, n12242, n12261, n12267, n12268,
         n12269, n12271, n12272, n12291, n12297, n12298, n12299, n12320,
         n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12332,
         n12334, n12336, n12338, n12340, n12342, n12344, n12346, n12348,
         n12351, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
         n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371,
         n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379,
         n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387,
         n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395,
         n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403,
         n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411,
         n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419,
         n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427,
         n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435,
         n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443,
         n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451,
         n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459,
         n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
         n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
         n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
         n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
         n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
         n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
         n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
         n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
         n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
         n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
         n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
         n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
         n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
         n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
         n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
         n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
         n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
         n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
         n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
         n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
         n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
         n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
         n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683,
         n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
         n12692, n12693, n12694, n12696, n12697, n12698, n12699, n12700,
         n12701, n12702, n12704, n12705, n12706, n12707, n12708, n12709,
         n12710, n12711, n12712, n12713, n12714, n12716, n12717, n12718,
         n12719, n12720, n12721, n12722, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12756, n12757, n12758, n12759, n12760, n12761, n12762,
         n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771,
         n12772, n12774, n12775, n12776, n12777, n12778, n12779, n12780,
         n12781, n12782, n12784, n12785, n12786, n12787, n12788, n12794,
         n12802, n12803, n12804, n12805, n12806, n12808, n12809, n12810,
         n12811, n12812, n12813, n12815, n12816, n12820, n12821, n12822,
         n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830,
         n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838,
         n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846,
         n12847, n12849, n12851, n12853, n12855, n12857, n12859, n12861,
         n12863, n12865, n12867, n12870, n12871, n12872, n12873, n12874,
         n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882,
         n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890,
         n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,
         n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906,
         n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
         n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922,
         n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930,
         n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938,
         n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946,
         n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954,
         n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962,
         n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970,
         n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978,
         n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986,
         n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994,
         n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002,
         n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010,
         n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
         n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026,
         n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
         n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042,
         n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,
         n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058,
         n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,
         n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074,
         n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082,
         n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090,
         n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098,
         n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
         n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114,
         n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122,
         n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130,
         n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
         n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146,
         n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,
         n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
         n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170,
         n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
         n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,
         n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194,
         n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
         n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
         n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218,
         n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,
         n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234,
         n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242,
         n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250,
         n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
         n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266,
         n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
         n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282,
         n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290,
         n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
         n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
         n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314,
         n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322,
         n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
         n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338,
         n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,
         n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
         n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362,
         n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
         n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
         n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
         n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394,
         n13395, n13396, n13397, n13398, n13399, n13401, n13412, n13435,
         n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443,
         n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451,
         n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459,
         n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ,
         \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ,
         \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ,
         \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ,
         \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ,
         \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ,
         \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ,
         \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ,
         \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ,
         \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ,
         \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ,
         \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ,
         \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ,
         \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ,
         \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ,
         \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ,
         \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ,
         \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ,
         \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ,
         \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ,
         \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ,
         \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ,
         \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ,
         \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ,
         \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ,
         \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ,
         \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ,
         \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ,
         \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ,
         \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ,
         \fadd_0_0_0_0_9/add_859/B[1] , \fadd_0_0_0_0_9/sub_784/B[0] ,
         \fadd_0_0_0_0_9/sub_784/B[1] , \fadd_0_0_0_0_8/add_859/B[1] ,
         \fadd_0_0_0_0_8/sub_784/B[0] , \fadd_0_0_0_0_8/sub_784/B[1] ,
         \fadd_0_0_0_0_7/add_859/B[1] , \fadd_0_0_0_0_7/sub_784/B[0] ,
         \fadd_0_0_0_0_7/sub_784/B[1] , \fadd_0_0_0_0_6/add_859/B[1] ,
         \fadd_0_0_0_0_6/sub_784/B[0] , \fadd_0_0_0_0_6/sub_784/B[1] ,
         \fadd_0_0_0_0_5/add_859/B[1] , \fadd_0_0_0_0_5/sub_784/B[0] ,
         \fadd_0_0_0_0_5/sub_784/B[1] , \fadd_0_0_0_0_4/add_859/B[1] ,
         \fadd_0_0_0_0_4/sub_784/B[0] , \fadd_0_0_0_0_4/sub_784/B[1] ,
         \fadd_0_0_0_0_3/add_859/B[1] , \fadd_0_0_0_0_3/sub_784/B[0] ,
         \fadd_0_0_0_0_3/sub_784/B[1] , \fadd_0_0_0_0_2/add_859/B[1] ,
         \fadd_0_0_0_0_2/sub_784/B[0] , \fadd_0_0_0_0_2/sub_784/B[1] ,
         \fadd_0_0_0_0_1/add_859/B[1] , \fadd_0_0_0_0_1/sub_784/B[0] ,
         \fadd_0_0_0_0_1/sub_784/B[1] , \fadd_0_0_0_0_0/add_859/B[1] ,
         \fadd_0_0_0_0_0/sub_784/B[0] , \fadd_0_0_0_0_0/sub_784/B[1] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/B[0] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/B[1] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/A[0] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/A[1] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/A[2] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/A[3] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/A[4] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/A[5] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/B[0] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/B[1] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/A[0] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/A[1] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/A[2] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/A[3] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/A[4] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/A[5] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/B[0] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/B[1] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/A[0] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/A[1] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/A[2] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/A[3] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/A[4] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/A[5] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/B[0] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/B[1] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/A[0] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/A[1] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/A[2] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/A[3] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/A[4] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/A[5] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/B[0] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/B[1] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/A[0] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/A[1] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/A[2] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/A[3] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/A[4] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/A[5] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/B[0] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/B[1] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/A[0] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/A[1] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/A[2] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/A[3] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/A[4] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/A[5] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/B[0] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/B[1] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/A[0] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/A[1] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/A[2] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/A[3] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/A[4] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/A[5] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/B[0] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/B[1] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/A[0] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/A[1] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/A[2] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/A[3] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/A[4] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/A[5] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/B[0] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/B[1] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/A[0] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/A[1] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/A[2] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/A[3] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/A[4] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/A[5] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/B[0] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/B[1] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/A[0] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/A[1] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/A[2] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/A[3] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/A[4] ,
         \add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/A[5] ,
         \add_0_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ,
         \add_0_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[2] ,
         \add_0_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[3] ,
         \add_0_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[4] ,
         \add_0_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[5] ,
         \sub_2_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[3] ,
         \sub_2_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[4] ,
         \add_0_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ,
         \add_0_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[2] ,
         \add_0_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[3] ,
         \add_0_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[4] ,
         \add_0_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[5] ,
         \sub_2_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[3] ,
         \sub_2_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[4] ,
         \add_0_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ,
         \add_0_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[2] ,
         \add_0_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[3] ,
         \add_0_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[4] ,
         \add_0_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[5] ,
         \sub_2_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[3] ,
         \sub_2_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[4] ,
         \add_0_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ,
         \add_0_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[2] ,
         \add_0_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[3] ,
         \add_0_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[4] ,
         \add_0_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[5] ,
         \sub_2_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[3] ,
         \sub_2_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[4] ,
         \add_0_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ,
         \add_0_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[2] ,
         \add_0_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[3] ,
         \add_0_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[4] ,
         \add_0_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[5] ,
         \sub_2_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[3] ,
         \sub_2_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[4] ,
         \add_0_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ,
         \add_0_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[2] ,
         \add_0_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[3] ,
         \add_0_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[4] ,
         \add_0_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[5] ,
         \sub_2_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[3] ,
         \sub_2_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[4] ,
         \add_0_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ,
         \add_0_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[2] ,
         \add_0_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[3] ,
         \add_0_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[4] ,
         \add_0_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[5] ,
         \sub_2_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[3] ,
         \sub_2_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[4] ,
         \add_0_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ,
         \add_0_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[2] ,
         \add_0_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[3] ,
         \add_0_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[4] ,
         \add_0_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[5] ,
         \sub_2_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[3] ,
         \sub_2_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[4] ,
         \add_0_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ,
         \add_0_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[2] ,
         \add_0_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[3] ,
         \add_0_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[4] ,
         \add_0_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[5] ,
         \sub_2_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[3] ,
         \sub_2_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[4] ,
         \add_0_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ,
         \add_0_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[2] ,
         \add_0_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[3] ,
         \add_0_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[4] ,
         \add_0_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[5] ,
         \sub_2_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[3] ,
         \sub_2_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[4] ,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
         n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
         n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722,
         n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
         n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
         n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,
         n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,
         n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
         n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,
         n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
         n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
         n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226,
         n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,
         n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
         n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,
         n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
         n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
         n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
         n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,
         n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
         n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298,
         n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,
         n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314,
         n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322,
         n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330,
         n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338,
         n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346,
         n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354,
         n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,
         n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370,
         n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378,
         n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386,
         n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394,
         n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402,
         n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410,
         n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418,
         n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426,
         n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434,
         n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442,
         n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450,
         n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458,
         n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466,
         n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474,
         n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482,
         n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490,
         n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
         n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,
         n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514,
         n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,
         n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,
         n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538,
         n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,
         n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
         n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562,
         n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
         n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
         n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586,
         n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,
         n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602,
         n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,
         n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
         n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,
         n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634,
         n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
         n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
         n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658,
         n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666,
         n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674,
         n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682,
         n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,
         n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
         n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706,
         n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
         n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,
         n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730,
         n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738,
         n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746,
         n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754,
         n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762,
         n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
         n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778,
         n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,
         n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794,
         n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802,
         n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810,
         n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818,
         n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826,
         n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834,
         n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
         n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850,
         n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
         n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
         n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,
         n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
         n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890,
         n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898,
         n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906,
         n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
         n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,
         n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
         n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938,
         n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946,
         n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
         n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962,
         n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970,
         n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978,
         n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,
         n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
         n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002;
  wire   [3:0] \fadd_0_0_0_0_0/syncexnxy_d1 ;
  wire   [9:0] \fadd_0_0_0_0_0/syncx_d2 ;
  wire   [9:0] \fadd_0_0_0_0_0/syncx_d1 ;
  wire   [10:0] \fadd_0_0_0_0_0/resultrounded ;
  wire   [10:0] \fadd_0_0_0_0_0/resultbeforeround ;
  wire   [6:0] \fadd_0_0_0_0_0/exponentresultfar1 ;
  wire   [6:0] \fadd_0_0_0_0_0/exponentresultfar0_d2 ;
  wire   [6:0] \fadd_0_0_0_0_0/exponentresultfar0_d1 ;
  wire   [7:0] \fadd_0_0_0_0_0/fracresultfar0 ;
  wire   [7:0] \fadd_0_0_0_0_0/fracyfarxorop ;
  wire   [6:0] \fadd_0_0_0_0_0/exponentresultclose_d1 ;
  wire   [4:0] \fadd_0_0_0_0_0/exponentresultclose ;
  wire   [5:0] \fadd_0_0_0_0_0/fracrclose1 ;
  wire   [6:0] \fadd_0_0_0_0_0/fracrcloseymx ;
  wire   [6:0] \fadd_0_0_0_0_0/fracrclosexmy ;
  wire   [5:0] \fadd_0_0_0_0_0/fracyclose1 ;
  wire   [8:4] \fadd_0_0_0_0_0/newx_d1 ;
  wire   [11:0] \fadd_0_0_0_0_0/newx ;
  wire   [4:0] \fadd_0_0_0_0_0/exponentdifferenceyx ;
  wire   [5:0] \fadd_0_0_0_0_0/exponentdifferencexy ;
  wire   [3:0] \fadd_0_0_0_0_1/syncexnxy_d1 ;
  wire   [9:0] \fadd_0_0_0_0_1/syncx_d2 ;
  wire   [9:0] \fadd_0_0_0_0_1/syncx_d1 ;
  wire   [10:0] \fadd_0_0_0_0_1/resultrounded ;
  wire   [10:0] \fadd_0_0_0_0_1/resultbeforeround ;
  wire   [6:0] \fadd_0_0_0_0_1/exponentresultfar1 ;
  wire   [6:0] \fadd_0_0_0_0_1/exponentresultfar0_d2 ;
  wire   [6:0] \fadd_0_0_0_0_1/exponentresultfar0_d1 ;
  wire   [7:0] \fadd_0_0_0_0_1/fracresultfar0 ;
  wire   [7:0] \fadd_0_0_0_0_1/fracyfarxorop ;
  wire   [6:0] \fadd_0_0_0_0_1/exponentresultclose_d1 ;
  wire   [4:0] \fadd_0_0_0_0_1/exponentresultclose ;
  wire   [5:0] \fadd_0_0_0_0_1/fracrclose1 ;
  wire   [6:0] \fadd_0_0_0_0_1/fracrcloseymx ;
  wire   [6:0] \fadd_0_0_0_0_1/fracrclosexmy ;
  wire   [5:0] \fadd_0_0_0_0_1/fracyclose1 ;
  wire   [8:4] \fadd_0_0_0_0_1/newx_d1 ;
  wire   [11:0] \fadd_0_0_0_0_1/newx ;
  wire   [4:0] \fadd_0_0_0_0_1/exponentdifferenceyx ;
  wire   [5:0] \fadd_0_0_0_0_1/exponentdifferencexy ;
  wire   [3:0] \fadd_0_0_0_0_2/syncexnxy_d1 ;
  wire   [9:0] \fadd_0_0_0_0_2/syncx_d2 ;
  wire   [9:0] \fadd_0_0_0_0_2/syncx_d1 ;
  wire   [10:0] \fadd_0_0_0_0_2/resultrounded ;
  wire   [10:0] \fadd_0_0_0_0_2/resultbeforeround ;
  wire   [6:0] \fadd_0_0_0_0_2/exponentresultfar1 ;
  wire   [6:0] \fadd_0_0_0_0_2/exponentresultfar0_d2 ;
  wire   [6:0] \fadd_0_0_0_0_2/exponentresultfar0_d1 ;
  wire   [7:0] \fadd_0_0_0_0_2/fracresultfar0 ;
  wire   [7:0] \fadd_0_0_0_0_2/fracyfarxorop ;
  wire   [6:0] \fadd_0_0_0_0_2/exponentresultclose_d1 ;
  wire   [4:0] \fadd_0_0_0_0_2/exponentresultclose ;
  wire   [5:0] \fadd_0_0_0_0_2/fracrclose1 ;
  wire   [6:0] \fadd_0_0_0_0_2/fracrcloseymx ;
  wire   [6:0] \fadd_0_0_0_0_2/fracrclosexmy ;
  wire   [5:0] \fadd_0_0_0_0_2/fracyclose1 ;
  wire   [8:4] \fadd_0_0_0_0_2/newx_d1 ;
  wire   [11:0] \fadd_0_0_0_0_2/newx ;
  wire   [4:0] \fadd_0_0_0_0_2/exponentdifferenceyx ;
  wire   [5:0] \fadd_0_0_0_0_2/exponentdifferencexy ;
  wire   [3:0] \fadd_0_0_0_0_3/syncexnxy_d1 ;
  wire   [9:0] \fadd_0_0_0_0_3/syncx_d2 ;
  wire   [9:0] \fadd_0_0_0_0_3/syncx_d1 ;
  wire   [10:0] \fadd_0_0_0_0_3/resultrounded ;
  wire   [10:0] \fadd_0_0_0_0_3/resultbeforeround ;
  wire   [6:0] \fadd_0_0_0_0_3/exponentresultfar1 ;
  wire   [6:0] \fadd_0_0_0_0_3/exponentresultfar0_d2 ;
  wire   [6:0] \fadd_0_0_0_0_3/exponentresultfar0_d1 ;
  wire   [7:0] \fadd_0_0_0_0_3/fracresultfar0 ;
  wire   [7:0] \fadd_0_0_0_0_3/fracyfarxorop ;
  wire   [6:0] \fadd_0_0_0_0_3/exponentresultclose_d1 ;
  wire   [4:0] \fadd_0_0_0_0_3/exponentresultclose ;
  wire   [5:0] \fadd_0_0_0_0_3/fracrclose1 ;
  wire   [6:0] \fadd_0_0_0_0_3/fracrcloseymx ;
  wire   [6:0] \fadd_0_0_0_0_3/fracrclosexmy ;
  wire   [5:0] \fadd_0_0_0_0_3/fracyclose1 ;
  wire   [8:4] \fadd_0_0_0_0_3/newx_d1 ;
  wire   [11:0] \fadd_0_0_0_0_3/newx ;
  wire   [4:0] \fadd_0_0_0_0_3/exponentdifferenceyx ;
  wire   [5:0] \fadd_0_0_0_0_3/exponentdifferencexy ;
  wire   [3:0] \fadd_0_0_0_0_4/syncexnxy_d1 ;
  wire   [9:0] \fadd_0_0_0_0_4/syncx_d2 ;
  wire   [9:0] \fadd_0_0_0_0_4/syncx_d1 ;
  wire   [10:0] \fadd_0_0_0_0_4/resultrounded ;
  wire   [10:0] \fadd_0_0_0_0_4/resultbeforeround ;
  wire   [6:0] \fadd_0_0_0_0_4/exponentresultfar1 ;
  wire   [6:0] \fadd_0_0_0_0_4/exponentresultfar0_d2 ;
  wire   [6:0] \fadd_0_0_0_0_4/exponentresultfar0_d1 ;
  wire   [7:0] \fadd_0_0_0_0_4/fracresultfar0 ;
  wire   [7:0] \fadd_0_0_0_0_4/fracyfarxorop ;
  wire   [6:0] \fadd_0_0_0_0_4/exponentresultclose_d1 ;
  wire   [4:0] \fadd_0_0_0_0_4/exponentresultclose ;
  wire   [5:0] \fadd_0_0_0_0_4/fracrclose1 ;
  wire   [6:0] \fadd_0_0_0_0_4/fracrcloseymx ;
  wire   [6:0] \fadd_0_0_0_0_4/fracrclosexmy ;
  wire   [5:0] \fadd_0_0_0_0_4/fracyclose1 ;
  wire   [8:4] \fadd_0_0_0_0_4/newx_d1 ;
  wire   [11:0] \fadd_0_0_0_0_4/newx ;
  wire   [4:0] \fadd_0_0_0_0_4/exponentdifferenceyx ;
  wire   [5:0] \fadd_0_0_0_0_4/exponentdifferencexy ;
  wire   [3:0] \fadd_0_0_0_0_5/syncexnxy_d1 ;
  wire   [9:0] \fadd_0_0_0_0_5/syncx_d2 ;
  wire   [9:0] \fadd_0_0_0_0_5/syncx_d1 ;
  wire   [10:0] \fadd_0_0_0_0_5/resultrounded ;
  wire   [10:0] \fadd_0_0_0_0_5/resultbeforeround ;
  wire   [6:0] \fadd_0_0_0_0_5/exponentresultfar1 ;
  wire   [6:0] \fadd_0_0_0_0_5/exponentresultfar0_d2 ;
  wire   [6:0] \fadd_0_0_0_0_5/exponentresultfar0_d1 ;
  wire   [7:0] \fadd_0_0_0_0_5/fracresultfar0 ;
  wire   [7:0] \fadd_0_0_0_0_5/fracyfarxorop ;
  wire   [6:0] \fadd_0_0_0_0_5/exponentresultclose_d1 ;
  wire   [4:0] \fadd_0_0_0_0_5/exponentresultclose ;
  wire   [5:0] \fadd_0_0_0_0_5/fracrclose1 ;
  wire   [6:0] \fadd_0_0_0_0_5/fracrcloseymx ;
  wire   [6:0] \fadd_0_0_0_0_5/fracrclosexmy ;
  wire   [5:0] \fadd_0_0_0_0_5/fracyclose1 ;
  wire   [8:4] \fadd_0_0_0_0_5/newx_d1 ;
  wire   [11:0] \fadd_0_0_0_0_5/newx ;
  wire   [4:0] \fadd_0_0_0_0_5/exponentdifferenceyx ;
  wire   [5:0] \fadd_0_0_0_0_5/exponentdifferencexy ;
  wire   [3:0] \fadd_0_0_0_0_6/syncexnxy_d1 ;
  wire   [9:0] \fadd_0_0_0_0_6/syncx_d2 ;
  wire   [9:0] \fadd_0_0_0_0_6/syncx_d1 ;
  wire   [10:0] \fadd_0_0_0_0_6/resultrounded ;
  wire   [10:0] \fadd_0_0_0_0_6/resultbeforeround ;
  wire   [6:0] \fadd_0_0_0_0_6/exponentresultfar1 ;
  wire   [6:0] \fadd_0_0_0_0_6/exponentresultfar0_d2 ;
  wire   [6:0] \fadd_0_0_0_0_6/exponentresultfar0_d1 ;
  wire   [7:0] \fadd_0_0_0_0_6/fracresultfar0 ;
  wire   [7:0] \fadd_0_0_0_0_6/fracyfarxorop ;
  wire   [6:0] \fadd_0_0_0_0_6/exponentresultclose_d1 ;
  wire   [4:0] \fadd_0_0_0_0_6/exponentresultclose ;
  wire   [5:0] \fadd_0_0_0_0_6/fracrclose1 ;
  wire   [6:0] \fadd_0_0_0_0_6/fracrcloseymx ;
  wire   [6:0] \fadd_0_0_0_0_6/fracrclosexmy ;
  wire   [5:0] \fadd_0_0_0_0_6/fracyclose1 ;
  wire   [8:4] \fadd_0_0_0_0_6/newx_d1 ;
  wire   [11:0] \fadd_0_0_0_0_6/newx ;
  wire   [4:0] \fadd_0_0_0_0_6/exponentdifferenceyx ;
  wire   [5:0] \fadd_0_0_0_0_6/exponentdifferencexy ;
  wire   [3:0] \fadd_0_0_0_0_7/syncexnxy_d1 ;
  wire   [9:0] \fadd_0_0_0_0_7/syncx_d2 ;
  wire   [9:0] \fadd_0_0_0_0_7/syncx_d1 ;
  wire   [10:0] \fadd_0_0_0_0_7/resultrounded ;
  wire   [10:0] \fadd_0_0_0_0_7/resultbeforeround ;
  wire   [6:0] \fadd_0_0_0_0_7/exponentresultfar1 ;
  wire   [6:0] \fadd_0_0_0_0_7/exponentresultfar0_d2 ;
  wire   [6:0] \fadd_0_0_0_0_7/exponentresultfar0_d1 ;
  wire   [7:0] \fadd_0_0_0_0_7/fracresultfar0 ;
  wire   [7:0] \fadd_0_0_0_0_7/fracyfarxorop ;
  wire   [6:0] \fadd_0_0_0_0_7/exponentresultclose_d1 ;
  wire   [4:0] \fadd_0_0_0_0_7/exponentresultclose ;
  wire   [5:0] \fadd_0_0_0_0_7/fracrclose1 ;
  wire   [6:0] \fadd_0_0_0_0_7/fracrcloseymx ;
  wire   [6:0] \fadd_0_0_0_0_7/fracrclosexmy ;
  wire   [5:0] \fadd_0_0_0_0_7/fracyclose1 ;
  wire   [8:4] \fadd_0_0_0_0_7/newx_d1 ;
  wire   [11:0] \fadd_0_0_0_0_7/newx ;
  wire   [4:0] \fadd_0_0_0_0_7/exponentdifferenceyx ;
  wire   [5:0] \fadd_0_0_0_0_7/exponentdifferencexy ;
  wire   [3:0] \fadd_0_0_0_0_8/syncexnxy_d1 ;
  wire   [9:0] \fadd_0_0_0_0_8/syncx_d2 ;
  wire   [9:0] \fadd_0_0_0_0_8/syncx_d1 ;
  wire   [10:0] \fadd_0_0_0_0_8/resultrounded ;
  wire   [10:0] \fadd_0_0_0_0_8/resultbeforeround ;
  wire   [6:0] \fadd_0_0_0_0_8/exponentresultfar1 ;
  wire   [6:0] \fadd_0_0_0_0_8/exponentresultfar0_d2 ;
  wire   [6:0] \fadd_0_0_0_0_8/exponentresultfar0_d1 ;
  wire   [7:0] \fadd_0_0_0_0_8/fracresultfar0 ;
  wire   [7:0] \fadd_0_0_0_0_8/fracyfarxorop ;
  wire   [6:0] \fadd_0_0_0_0_8/exponentresultclose_d1 ;
  wire   [4:0] \fadd_0_0_0_0_8/exponentresultclose ;
  wire   [5:0] \fadd_0_0_0_0_8/fracrclose1 ;
  wire   [6:0] \fadd_0_0_0_0_8/fracrcloseymx ;
  wire   [6:0] \fadd_0_0_0_0_8/fracrclosexmy ;
  wire   [5:0] \fadd_0_0_0_0_8/fracyclose1 ;
  wire   [8:4] \fadd_0_0_0_0_8/newx_d1 ;
  wire   [11:0] \fadd_0_0_0_0_8/newx ;
  wire   [4:0] \fadd_0_0_0_0_8/exponentdifferenceyx ;
  wire   [5:0] \fadd_0_0_0_0_8/exponentdifferencexy ;
  wire   [3:0] \fadd_0_0_0_0_9/syncexnxy_d1 ;
  wire   [9:0] \fadd_0_0_0_0_9/syncx_d2 ;
  wire   [9:0] \fadd_0_0_0_0_9/syncx_d1 ;
  wire   [10:0] \fadd_0_0_0_0_9/resultrounded ;
  wire   [10:0] \fadd_0_0_0_0_9/resultbeforeround ;
  wire   [6:0] \fadd_0_0_0_0_9/exponentresultfar1 ;
  wire   [6:0] \fadd_0_0_0_0_9/exponentresultfar0_d2 ;
  wire   [6:0] \fadd_0_0_0_0_9/exponentresultfar0_d1 ;
  wire   [7:0] \fadd_0_0_0_0_9/fracresultfar0 ;
  wire   [7:0] \fadd_0_0_0_0_9/fracyfarxorop ;
  wire   [6:0] \fadd_0_0_0_0_9/exponentresultclose_d1 ;
  wire   [4:0] \fadd_0_0_0_0_9/exponentresultclose ;
  wire   [5:0] \fadd_0_0_0_0_9/fracrclose1 ;
  wire   [6:0] \fadd_0_0_0_0_9/fracrcloseymx ;
  wire   [6:0] \fadd_0_0_0_0_9/fracrclosexmy ;
  wire   [5:0] \fadd_0_0_0_0_9/fracyclose1 ;
  wire   [8:4] \fadd_0_0_0_0_9/newx_d1 ;
  wire   [11:0] \fadd_0_0_0_0_9/newx ;
  wire   [4:0] \fadd_0_0_0_0_9/exponentdifferenceyx ;
  wire   [5:0] \fadd_0_0_0_0_9/exponentdifferencexy ;
  wire   [5:0] \fadd_0_0_0_0_0/norm/level1 ;
  wire   [5:0] \fadd_0_0_0_0_1/norm/level1 ;
  wire   [5:0] \fadd_0_0_0_0_2/norm/level1 ;
  wire   [5:0] \fadd_0_0_0_0_3/norm/level1 ;
  wire   [5:0] \fadd_0_0_0_0_4/norm/level1 ;
  wire   [5:0] \fadd_0_0_0_0_5/norm/level1 ;
  wire   [5:0] \fadd_0_0_0_0_6/norm/level1 ;
  wire   [5:0] \fadd_0_0_0_0_7/norm/level1 ;
  wire   [5:0] \fadd_0_0_0_0_8/norm/level1 ;
  wire   [5:0] \fadd_0_0_0_0_9/norm/level1 ;
  wire   [2:0] \fadd_0_0_0_0_0/rightshiftercomponent/ps_d1 ;
  wire   [2:0] \fadd_0_0_0_0_1/rightshiftercomponent/ps_d1 ;
  wire   [2:0] \fadd_0_0_0_0_2/rightshiftercomponent/ps_d1 ;
  wire   [2:0] \fadd_0_0_0_0_3/rightshiftercomponent/ps_d1 ;
  wire   [2:0] \fadd_0_0_0_0_4/rightshiftercomponent/ps_d1 ;
  wire   [2:0] \fadd_0_0_0_0_5/rightshiftercomponent/ps_d1 ;
  wire   [2:0] \fadd_0_0_0_0_6/rightshiftercomponent/ps_d1 ;
  wire   [2:0] \fadd_0_0_0_0_7/rightshiftercomponent/ps_d1 ;
  wire   [2:0] \fadd_0_0_0_0_8/rightshiftercomponent/ps_d1 ;
  wire   [2:0] \fadd_0_0_0_0_9/rightshiftercomponent/ps_d1 ;
  wire   [7:0] \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/y_d2 ;
  wire   [7:0] \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/y_d1 ;
  wire   [7:0] \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/x_d2 ;
  wire   [7:0] \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/x_d1 ;
  wire   [7:0] \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/y_d2 ;
  wire   [7:0] \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/y_d1 ;
  wire   [7:0] \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/x_d2 ;
  wire   [7:0] \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/x_d1 ;
  wire   [7:0] \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/y_d2 ;
  wire   [7:0] \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/y_d1 ;
  wire   [7:0] \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/x_d2 ;
  wire   [7:0] \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/x_d1 ;
  wire   [7:0] \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/y_d2 ;
  wire   [7:0] \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/y_d1 ;
  wire   [7:0] \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/x_d2 ;
  wire   [7:0] \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/x_d1 ;
  wire   [7:0] \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/y_d2 ;
  wire   [7:0] \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/y_d1 ;
  wire   [7:0] \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/x_d2 ;
  wire   [7:0] \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/x_d1 ;
  wire   [7:0] \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/y_d2 ;
  wire   [7:0] \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/y_d1 ;
  wire   [7:0] \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/x_d2 ;
  wire   [7:0] \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/x_d1 ;
  wire   [7:0] \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/y_d2 ;
  wire   [7:0] \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/y_d1 ;
  wire   [7:0] \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/x_d2 ;
  wire   [7:0] \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/x_d1 ;
  wire   [7:0] \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/y_d2 ;
  wire   [7:0] \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/y_d1 ;
  wire   [7:0] \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/x_d2 ;
  wire   [7:0] \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/x_d1 ;
  wire   [7:0] \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/y_d2 ;
  wire   [7:0] \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/y_d1 ;
  wire   [7:0] \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/x_d2 ;
  wire   [7:0] \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/x_d1 ;
  wire   [7:0] \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/y_d2 ;
  wire   [7:0] \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/y_d1 ;
  wire   [7:0] \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/x_d2 ;
  wire   [7:0] \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/x_d1 ;
  wire   [7:0] \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/y_d1 ;
  wire   [7:0] \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/x_d1 ;
  wire   [10:9] \fmul_0_0_0_0_0/expsigpostround ;
  wire   [9:1] \fmul_0_0_0_0_0/sigprodext ;
  wire   [6:0] \fmul_0_0_0_0_0/exppostnorm ;
  wire   [1:0] \fmul_0_0_0_0_0/exc ;
  wire   [9:0] \fmul_0_0_0_0_0/sigprod ;
  wire   [10:9] \fmul_0_0_0_0_1/expsigpostround ;
  wire   [9:1] \fmul_0_0_0_0_1/sigprodext ;
  wire   [6:0] \fmul_0_0_0_0_1/exppostnorm ;
  wire   [1:0] \fmul_0_0_0_0_1/exc ;
  wire   [9:0] \fmul_0_0_0_0_1/sigprod ;
  wire   [10:9] \fmul_0_0_0_0_2/expsigpostround ;
  wire   [9:1] \fmul_0_0_0_0_2/sigprodext ;
  wire   [6:0] \fmul_0_0_0_0_2/exppostnorm ;
  wire   [1:0] \fmul_0_0_0_0_2/exc ;
  wire   [9:0] \fmul_0_0_0_0_2/sigprod ;
  wire   [10:9] \fmul_0_0_0_0_3/expsigpostround ;
  wire   [9:1] \fmul_0_0_0_0_3/sigprodext ;
  wire   [6:0] \fmul_0_0_0_0_3/exppostnorm ;
  wire   [1:0] \fmul_0_0_0_0_3/exc ;
  wire   [9:0] \fmul_0_0_0_0_3/sigprod ;
  wire   [10:9] \fmul_0_0_0_0_4/expsigpostround ;
  wire   [9:1] \fmul_0_0_0_0_4/sigprodext ;
  wire   [6:0] \fmul_0_0_0_0_4/exppostnorm ;
  wire   [1:0] \fmul_0_0_0_0_4/exc ;
  wire   [9:0] \fmul_0_0_0_0_4/sigprod ;
  wire   [10:9] \fmul_0_0_0_0_5/expsigpostround ;
  wire   [9:1] \fmul_0_0_0_0_5/sigprodext ;
  wire   [6:0] \fmul_0_0_0_0_5/exppostnorm ;
  wire   [1:0] \fmul_0_0_0_0_5/exc ;
  wire   [9:0] \fmul_0_0_0_0_5/sigprod ;
  wire   [10:9] \fmul_0_0_0_0_6/expsigpostround ;
  wire   [9:1] \fmul_0_0_0_0_6/sigprodext ;
  wire   [6:0] \fmul_0_0_0_0_6/exppostnorm ;
  wire   [1:0] \fmul_0_0_0_0_6/exc ;
  wire   [9:0] \fmul_0_0_0_0_6/sigprod ;
  wire   [10:9] \fmul_0_0_0_0_7/expsigpostround ;
  wire   [9:1] \fmul_0_0_0_0_7/sigprodext ;
  wire   [6:0] \fmul_0_0_0_0_7/exppostnorm ;
  wire   [1:0] \fmul_0_0_0_0_7/exc ;
  wire   [9:0] \fmul_0_0_0_0_7/sigprod ;
  wire   [9:1] \fmul_0_0_0_0_8/sigprodext ;
  wire   [6:0] \fmul_0_0_0_0_8/exppostnorm ;
  wire   [1:0] \fmul_0_0_0_0_8/exc ;
  wire   [9:0] \fmul_0_0_0_0_8/sigprod ;
  wire   [10:9] \fmul_0_0_0_0_9/expsigpostround ;
  wire   [9:1] \fmul_0_0_0_0_9/sigprodext ;
  wire   [6:0] \fmul_0_0_0_0_9/exppostnorm ;
  wire   [1:0] \fmul_0_0_0_0_9/exc ;
  wire   [9:0] \fmul_0_0_0_0_9/sigprod ;
  wire   [10:0] \fmul_0_0_0_0_0/roundingadder/x_1_d1 ;
  wire   [10:0] \fmul_0_0_0_0_1/roundingadder/x_1_d1 ;
  wire   [10:0] \fmul_0_0_0_0_2/roundingadder/x_1_d1 ;
  wire   [10:0] \fmul_0_0_0_0_3/roundingadder/x_1_d1 ;
  wire   [10:0] \fmul_0_0_0_0_4/roundingadder/x_1_d1 ;
  wire   [10:0] \fmul_0_0_0_0_5/roundingadder/x_1_d1 ;
  wire   [10:0] \fmul_0_0_0_0_6/roundingadder/x_1_d1 ;
  wire   [10:0] \fmul_0_0_0_0_7/roundingadder/x_1_d1 ;
  wire   [10:0] \fmul_0_0_0_0_8/roundingadder/x_1_d1 ;
  wire   [10:0] \fmul_0_0_0_0_9/roundingadder/x_1_d1 ;
  wire   [10:1] \add_1_root_fmul_0_0_0_0_9/roundingadder/add_57/carry ;
  wire   [10:1] \add_1_root_fmul_0_0_0_0_8/roundingadder/add_57/carry ;
  wire   [10:1] \add_1_root_fmul_0_0_0_0_7/roundingadder/add_57/carry ;
  wire   [10:1] \add_1_root_fmul_0_0_0_0_6/roundingadder/add_57/carry ;
  wire   [10:1] \add_1_root_fmul_0_0_0_0_5/roundingadder/add_57/carry ;
  wire   [10:1] \add_1_root_fmul_0_0_0_0_4/roundingadder/add_57/carry ;
  wire   [10:1] \add_1_root_fmul_0_0_0_0_3/roundingadder/add_57/carry ;
  wire   [10:1] \add_1_root_fmul_0_0_0_0_2/roundingadder/add_57/carry ;
  wire   [10:1] \add_1_root_fmul_0_0_0_0_1/roundingadder/add_57/carry ;
  wire   [10:1] \add_1_root_fmul_0_0_0_0_0/roundingadder/add_57/carry ;
  wire  
         [10:1] \add_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry 
;
  wire  
         [10:1] \add_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry 
;
  wire  
         [10:1] \add_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry 
;
  wire  
         [10:1] \add_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry 
;
  wire  
         [10:1] \add_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry 
;
  wire  
         [10:1] \add_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry 
;
  wire  
         [10:1] \add_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry 
;
  wire  
         [10:1] \add_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry 
;
  wire  
         [10:1] \add_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry 
;
  wire  
         [10:1] \add_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry 
;
  wire   [6:1] \fadd_0_0_0_0_9/add_859/carry ;
  wire   [6:0] \fadd_0_0_0_0_9/sub_784/carry ;
  wire   [5:0] \fadd_0_0_0_0_9/sub_710/carry ;
  wire   [6:0] \fadd_0_0_0_0_9/sub_707/carry ;
  wire   [6:1] \fadd_0_0_0_0_8/add_859/carry ;
  wire   [6:0] \fadd_0_0_0_0_8/sub_784/carry ;
  wire   [5:0] \fadd_0_0_0_0_8/sub_710/carry ;
  wire   [6:0] \fadd_0_0_0_0_8/sub_707/carry ;
  wire   [6:1] \fadd_0_0_0_0_7/add_859/carry ;
  wire   [6:0] \fadd_0_0_0_0_7/sub_784/carry ;
  wire   [5:0] \fadd_0_0_0_0_7/sub_710/carry ;
  wire   [6:0] \fadd_0_0_0_0_7/sub_707/carry ;
  wire   [6:1] \fadd_0_0_0_0_6/add_859/carry ;
  wire   [6:0] \fadd_0_0_0_0_6/sub_784/carry ;
  wire   [5:0] \fadd_0_0_0_0_6/sub_710/carry ;
  wire   [6:0] \fadd_0_0_0_0_6/sub_707/carry ;
  wire   [6:1] \fadd_0_0_0_0_5/add_859/carry ;
  wire   [6:0] \fadd_0_0_0_0_5/sub_784/carry ;
  wire   [5:0] \fadd_0_0_0_0_5/sub_710/carry ;
  wire   [6:0] \fadd_0_0_0_0_5/sub_707/carry ;
  wire   [6:1] \fadd_0_0_0_0_4/add_859/carry ;
  wire   [6:0] \fadd_0_0_0_0_4/sub_784/carry ;
  wire   [5:0] \fadd_0_0_0_0_4/sub_710/carry ;
  wire   [6:0] \fadd_0_0_0_0_4/sub_707/carry ;
  wire   [6:1] \fadd_0_0_0_0_3/add_859/carry ;
  wire   [6:0] \fadd_0_0_0_0_3/sub_784/carry ;
  wire   [5:0] \fadd_0_0_0_0_3/sub_710/carry ;
  wire   [6:0] \fadd_0_0_0_0_3/sub_707/carry ;
  wire   [6:1] \fadd_0_0_0_0_2/add_859/carry ;
  wire   [6:0] \fadd_0_0_0_0_2/sub_784/carry ;
  wire   [5:0] \fadd_0_0_0_0_2/sub_710/carry ;
  wire   [6:0] \fadd_0_0_0_0_2/sub_707/carry ;
  wire   [6:1] \fadd_0_0_0_0_1/add_859/carry ;
  wire   [6:0] \fadd_0_0_0_0_1/sub_784/carry ;
  wire   [5:0] \fadd_0_0_0_0_1/sub_710/carry ;
  wire   [6:0] \fadd_0_0_0_0_1/sub_707/carry ;
  wire   [6:1] \fadd_0_0_0_0_0/add_859/carry ;
  wire   [6:0] \fadd_0_0_0_0_0/sub_784/carry ;
  wire   [5:0] \fadd_0_0_0_0_0/sub_710/carry ;
  wire   [6:0] \fadd_0_0_0_0_0/sub_707/carry ;
  wire   [6:1] \add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/carry ;
  wire   [6:1] \add_2_root_sub_1_root_fmul_0_0_0_0_0/add_321/carry ;
  wire   [6:1] \add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/carry ;
  wire   [6:1] \add_2_root_sub_1_root_fmul_0_0_0_0_1/add_321/carry ;
  wire   [6:1] \add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/carry ;
  wire   [6:1] \add_2_root_sub_1_root_fmul_0_0_0_0_2/add_321/carry ;
  wire   [6:1] \add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/carry ;
  wire   [6:1] \add_2_root_sub_1_root_fmul_0_0_0_0_3/add_321/carry ;
  wire   [6:1] \add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/carry ;
  wire   [6:1] \add_2_root_sub_1_root_fmul_0_0_0_0_4/add_321/carry ;
  wire   [6:1] \add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/carry ;
  wire   [6:1] \add_2_root_sub_1_root_fmul_0_0_0_0_5/add_321/carry ;
  wire   [6:1] \add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/carry ;
  wire   [6:1] \add_2_root_sub_1_root_fmul_0_0_0_0_6/add_321/carry ;
  wire   [6:1] \add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/carry ;
  wire   [6:1] \add_2_root_sub_1_root_fmul_0_0_0_0_7/add_321/carry ;
  wire   [6:1] \add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/carry ;
  wire   [6:1] \add_2_root_sub_1_root_fmul_0_0_0_0_8/add_321/carry ;
  wire   [6:1] \add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/carry ;
  wire   [6:1] \add_2_root_sub_1_root_fmul_0_0_0_0_9/add_321/carry ;
  wire  
         [7:0] \sub_0_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry 
;
  wire  
         [6:1] \add_0_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry 
;
  wire  
         [7:0] \sub_0_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry 
;
  wire  
         [6:1] \add_0_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry 
;
  wire  
         [7:0] \sub_0_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry 
;
  wire  
         [6:1] \add_0_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry 
;
  wire  
         [7:0] \sub_0_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry 
;
  wire  
         [6:1] \add_0_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry 
;
  wire  
         [7:0] \sub_0_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry 
;
  wire  
         [6:1] \add_0_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry 
;
  wire  
         [7:0] \sub_0_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry 
;
  wire  
         [6:1] \add_0_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry 
;
  wire  
         [7:0] \sub_0_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry 
;
  wire  
         [6:1] \add_0_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry 
;
  wire  
         [7:0] \sub_0_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry 
;
  wire  
         [6:1] \add_0_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry 
;
  wire  
         [7:0] \sub_0_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry 
;
  wire  
         [6:1] \add_0_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry 
;
  wire  
         [7:0] \sub_0_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry 
;
  wire  
         [6:1] \add_0_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry 
;
  assign \U616/DATA2_0  = p__arg0_0_0[0];
  assign \U616/DATA2_1  = p__arg0_0_0[1];
  assign \U616/DATA2_2  = p__arg0_0_0[2];
  assign \U616/DATA2_3  = p__arg0_0_0[3];
  assign \U616/DATA2_4  = p__arg0_0_0[4];
  assign \U616/DATA2_5  = p__arg0_0_0[5];
  assign \U616/DATA2_6  = p__arg0_0_0[6];
  assign \U616/DATA2_7  = p__arg0_0_0[7];
  assign \U616/DATA2_8  = p__arg0_0_0[8];
  assign \U616/DATA2_9  = p__arg0_0_0[9];
  assign \U616/DATA2_10  = p__arg0_0_0[10];
  assign \U616/DATA2_11  = p__arg0_0_0[11];
  assign \U616/DATA1_0  = p__arg0_0_1[0];
  assign \U616/DATA1_1  = p__arg0_0_1[1];
  assign \U616/DATA1_2  = p__arg0_0_1[2];
  assign \U616/DATA1_3  = p__arg0_0_1[3];
  assign \U616/DATA1_4  = p__arg0_0_1[4];
  assign \U616/DATA1_5  = p__arg0_0_1[5];
  assign \U616/DATA1_6  = p__arg0_0_1[6];
  assign \U616/DATA1_7  = p__arg0_0_1[7];
  assign \U616/DATA1_8  = p__arg0_0_1[8];
  assign \U616/DATA1_9  = p__arg0_0_1[9];
  assign \U616/DATA1_10  = p__arg0_0_1[10];
  assign \U616/DATA1_11  = p__arg0_0_1[11];
  assign \U615/DATA2_0  = p___constant_11x11xf32_0_0[0];
  assign \U615/DATA2_1  = p___constant_11x11xf32_0_0[1];
  assign \U615/DATA2_2  = p___constant_11x11xf32_0_0[2];
  assign \U615/DATA2_3  = p___constant_11x11xf32_0_0[3];
  assign \U615/DATA2_4  = p___constant_11x11xf32_0_0[4];
  assign \U615/DATA2_5  = p___constant_11x11xf32_0_0[5];
  assign \U615/DATA2_6  = p___constant_11x11xf32_0_0[6];
  assign \U615/DATA2_7  = p___constant_11x11xf32_0_0[7];
  assign \U615/DATA2_8  = p___constant_11x11xf32_0_0[8];
  assign \U615/DATA2_9  = p___constant_11x11xf32_0_0[9];
  assign \U615/DATA2_10  = p___constant_11x11xf32_0_0[10];
  assign \U615/DATA2_11  = p___constant_11x11xf32_0_0[11];
  assign \U615/DATA1_0  = p___constant_11x11xf32_0_1[0];
  assign \U615/DATA1_1  = p___constant_11x11xf32_0_1[1];
  assign \U615/DATA1_2  = p___constant_11x11xf32_0_1[2];
  assign \U615/DATA1_3  = p___constant_11x11xf32_0_1[3];
  assign \U615/DATA1_4  = p___constant_11x11xf32_0_1[4];
  assign \U615/DATA1_5  = p___constant_11x11xf32_0_1[5];
  assign \U615/DATA1_6  = p___constant_11x11xf32_0_1[6];
  assign \U615/DATA1_7  = p___constant_11x11xf32_0_1[7];
  assign \U615/DATA1_8  = p___constant_11x11xf32_0_1[8];
  assign \U615/DATA1_9  = p___constant_11x11xf32_0_1[9];
  assign \U615/DATA1_10  = p___constant_11x11xf32_0_1[10];
  assign \U615/DATA1_11  = p___constant_11x11xf32_0_1[11];
  assign \U611/DATA1_0  = p__arg0_0_2[0];
  assign \U611/DATA1_1  = p__arg0_0_2[1];
  assign \U611/DATA1_2  = p__arg0_0_2[2];
  assign \U611/DATA1_3  = p__arg0_0_2[3];
  assign \U611/DATA1_4  = p__arg0_0_2[4];
  assign \U611/DATA1_5  = p__arg0_0_2[5];
  assign \U611/DATA1_6  = p__arg0_0_2[6];
  assign \U611/DATA1_7  = p__arg0_0_2[7];
  assign \U611/DATA1_8  = p__arg0_0_2[8];
  assign \U611/DATA1_9  = p__arg0_0_2[9];
  assign \U611/DATA1_10  = p__arg0_0_2[10];
  assign \U611/DATA1_11  = p__arg0_0_2[11];
  assign \U610/DATA1_0  = p___constant_11x11xf32_0_2[0];
  assign \U610/DATA1_1  = p___constant_11x11xf32_0_2[1];
  assign \U610/DATA1_2  = p___constant_11x11xf32_0_2[2];
  assign \U610/DATA1_3  = p___constant_11x11xf32_0_2[3];
  assign \U610/DATA1_4  = p___constant_11x11xf32_0_2[4];
  assign \U610/DATA1_5  = p___constant_11x11xf32_0_2[5];
  assign \U610/DATA1_6  = p___constant_11x11xf32_0_2[6];
  assign \U610/DATA1_7  = p___constant_11x11xf32_0_2[7];
  assign \U610/DATA1_8  = p___constant_11x11xf32_0_2[8];
  assign \U610/DATA1_9  = p___constant_11x11xf32_0_2[9];
  assign \U610/DATA1_10  = p___constant_11x11xf32_0_2[10];
  assign \U610/DATA1_11  = p___constant_11x11xf32_0_2[11];
  assign \U606/DATA1_0  = p__arg0_0_3[0];
  assign \U606/DATA1_1  = p__arg0_0_3[1];
  assign \U606/DATA1_2  = p__arg0_0_3[2];
  assign \U606/DATA1_3  = p__arg0_0_3[3];
  assign \U606/DATA1_4  = p__arg0_0_3[4];
  assign \U606/DATA1_5  = p__arg0_0_3[5];
  assign \U606/DATA1_6  = p__arg0_0_3[6];
  assign \U606/DATA1_7  = p__arg0_0_3[7];
  assign \U606/DATA1_8  = p__arg0_0_3[8];
  assign \U606/DATA1_9  = p__arg0_0_3[9];
  assign \U606/DATA1_10  = p__arg0_0_3[10];
  assign \U606/DATA1_11  = p__arg0_0_3[11];
  assign \U605/DATA1_0  = p___constant_11x11xf32_0_3[0];
  assign \U605/DATA1_1  = p___constant_11x11xf32_0_3[1];
  assign \U605/DATA1_2  = p___constant_11x11xf32_0_3[2];
  assign \U605/DATA1_3  = p___constant_11x11xf32_0_3[3];
  assign \U605/DATA1_4  = p___constant_11x11xf32_0_3[4];
  assign \U605/DATA1_5  = p___constant_11x11xf32_0_3[5];
  assign \U605/DATA1_6  = p___constant_11x11xf32_0_3[6];
  assign \U605/DATA1_7  = p___constant_11x11xf32_0_3[7];
  assign \U605/DATA1_8  = p___constant_11x11xf32_0_3[8];
  assign \U605/DATA1_9  = p___constant_11x11xf32_0_3[9];
  assign \U605/DATA1_10  = p___constant_11x11xf32_0_3[10];
  assign \U605/DATA1_11  = p___constant_11x11xf32_0_3[11];
  assign \U601/DATA1_0  = p__arg0_0_4[0];
  assign \U601/DATA1_1  = p__arg0_0_4[1];
  assign \U601/DATA1_2  = p__arg0_0_4[2];
  assign \U601/DATA1_3  = p__arg0_0_4[3];
  assign \U601/DATA1_4  = p__arg0_0_4[4];
  assign \U601/DATA1_5  = p__arg0_0_4[5];
  assign \U601/DATA1_6  = p__arg0_0_4[6];
  assign \U601/DATA1_7  = p__arg0_0_4[7];
  assign \U601/DATA1_8  = p__arg0_0_4[8];
  assign \U601/DATA1_9  = p__arg0_0_4[9];
  assign \U601/DATA1_10  = p__arg0_0_4[10];
  assign \U601/DATA1_11  = p__arg0_0_4[11];
  assign \U600/DATA1_0  = p___constant_11x11xf32_0_4[0];
  assign \U600/DATA1_1  = p___constant_11x11xf32_0_4[1];
  assign \U600/DATA1_2  = p___constant_11x11xf32_0_4[2];
  assign \U600/DATA1_3  = p___constant_11x11xf32_0_4[3];
  assign \U600/DATA1_4  = p___constant_11x11xf32_0_4[4];
  assign \U600/DATA1_5  = p___constant_11x11xf32_0_4[5];
  assign \U600/DATA1_6  = p___constant_11x11xf32_0_4[6];
  assign \U600/DATA1_7  = p___constant_11x11xf32_0_4[7];
  assign \U600/DATA1_8  = p___constant_11x11xf32_0_4[8];
  assign \U600/DATA1_9  = p___constant_11x11xf32_0_4[9];
  assign \U600/DATA1_10  = p___constant_11x11xf32_0_4[10];
  assign \U600/DATA1_11  = p___constant_11x11xf32_0_4[11];
  assign \U596/DATA1_0  = p__arg0_0_5[0];
  assign \U596/DATA1_1  = p__arg0_0_5[1];
  assign \U596/DATA1_2  = p__arg0_0_5[2];
  assign \U596/DATA1_3  = p__arg0_0_5[3];
  assign \U596/DATA1_4  = p__arg0_0_5[4];
  assign \U596/DATA1_5  = p__arg0_0_5[5];
  assign \U596/DATA1_6  = p__arg0_0_5[6];
  assign \U596/DATA1_7  = p__arg0_0_5[7];
  assign \U596/DATA1_8  = p__arg0_0_5[8];
  assign \U596/DATA1_9  = p__arg0_0_5[9];
  assign \U596/DATA1_10  = p__arg0_0_5[10];
  assign \U596/DATA1_11  = p__arg0_0_5[11];
  assign \U595/DATA1_0  = p___constant_11x11xf32_0_5[0];
  assign \U595/DATA1_1  = p___constant_11x11xf32_0_5[1];
  assign \U595/DATA1_2  = p___constant_11x11xf32_0_5[2];
  assign \U595/DATA1_3  = p___constant_11x11xf32_0_5[3];
  assign \U595/DATA1_4  = p___constant_11x11xf32_0_5[4];
  assign \U595/DATA1_5  = p___constant_11x11xf32_0_5[5];
  assign \U595/DATA1_6  = p___constant_11x11xf32_0_5[6];
  assign \U595/DATA1_7  = p___constant_11x11xf32_0_5[7];
  assign \U595/DATA1_8  = p___constant_11x11xf32_0_5[8];
  assign \U595/DATA1_9  = p___constant_11x11xf32_0_5[9];
  assign \U595/DATA1_10  = p___constant_11x11xf32_0_5[10];
  assign \U595/DATA1_11  = p___constant_11x11xf32_0_5[11];
  assign \U591/DATA1_0  = p__arg0_0_6[0];
  assign \U591/DATA1_1  = p__arg0_0_6[1];
  assign \U591/DATA1_2  = p__arg0_0_6[2];
  assign \U591/DATA1_3  = p__arg0_0_6[3];
  assign \U591/DATA1_4  = p__arg0_0_6[4];
  assign \U591/DATA1_5  = p__arg0_0_6[5];
  assign \U591/DATA1_6  = p__arg0_0_6[6];
  assign \U591/DATA1_7  = p__arg0_0_6[7];
  assign \U591/DATA1_8  = p__arg0_0_6[8];
  assign \U591/DATA1_9  = p__arg0_0_6[9];
  assign \U591/DATA1_10  = p__arg0_0_6[10];
  assign \U591/DATA1_11  = p__arg0_0_6[11];
  assign \U590/DATA1_0  = p___constant_11x11xf32_0_6[0];
  assign \U590/DATA1_1  = p___constant_11x11xf32_0_6[1];
  assign \U590/DATA1_2  = p___constant_11x11xf32_0_6[2];
  assign \U590/DATA1_3  = p___constant_11x11xf32_0_6[3];
  assign \U590/DATA1_4  = p___constant_11x11xf32_0_6[4];
  assign \U590/DATA1_5  = p___constant_11x11xf32_0_6[5];
  assign \U590/DATA1_6  = p___constant_11x11xf32_0_6[6];
  assign \U590/DATA1_7  = p___constant_11x11xf32_0_6[7];
  assign \U590/DATA1_8  = p___constant_11x11xf32_0_6[8];
  assign \U590/DATA1_9  = p___constant_11x11xf32_0_6[9];
  assign \U590/DATA1_10  = p___constant_11x11xf32_0_6[10];
  assign \U590/DATA1_11  = p___constant_11x11xf32_0_6[11];
  assign \U586/DATA1_0  = p__arg0_0_7[0];
  assign \U586/DATA1_1  = p__arg0_0_7[1];
  assign \U586/DATA1_2  = p__arg0_0_7[2];
  assign \U586/DATA1_3  = p__arg0_0_7[3];
  assign \U586/DATA1_4  = p__arg0_0_7[4];
  assign \U586/DATA1_5  = p__arg0_0_7[5];
  assign \U586/DATA1_6  = p__arg0_0_7[6];
  assign \U586/DATA1_7  = p__arg0_0_7[7];
  assign \U586/DATA1_8  = p__arg0_0_7[8];
  assign \U586/DATA1_9  = p__arg0_0_7[9];
  assign \U586/DATA1_10  = p__arg0_0_7[10];
  assign \U586/DATA1_11  = p__arg0_0_7[11];
  assign \U585/DATA1_0  = p___constant_11x11xf32_0_7[0];
  assign \U585/DATA1_1  = p___constant_11x11xf32_0_7[1];
  assign \U585/DATA1_2  = p___constant_11x11xf32_0_7[2];
  assign \U585/DATA1_3  = p___constant_11x11xf32_0_7[3];
  assign \U585/DATA1_4  = p___constant_11x11xf32_0_7[4];
  assign \U585/DATA1_5  = p___constant_11x11xf32_0_7[5];
  assign \U585/DATA1_6  = p___constant_11x11xf32_0_7[6];
  assign \U585/DATA1_7  = p___constant_11x11xf32_0_7[7];
  assign \U585/DATA1_8  = p___constant_11x11xf32_0_7[8];
  assign \U585/DATA1_9  = p___constant_11x11xf32_0_7[9];
  assign \U585/DATA1_10  = p___constant_11x11xf32_0_7[10];
  assign \U585/DATA1_11  = p___constant_11x11xf32_0_7[11];
  assign \U581/DATA1_0  = p__arg0_0_8[0];
  assign \U581/DATA1_1  = p__arg0_0_8[1];
  assign \U581/DATA1_2  = p__arg0_0_8[2];
  assign \U581/DATA1_3  = p__arg0_0_8[3];
  assign \U581/DATA1_4  = p__arg0_0_8[4];
  assign \U581/DATA1_5  = p__arg0_0_8[5];
  assign \U581/DATA1_6  = p__arg0_0_8[6];
  assign \U581/DATA1_7  = p__arg0_0_8[7];
  assign \U581/DATA1_8  = p__arg0_0_8[8];
  assign \U581/DATA1_9  = p__arg0_0_8[9];
  assign \U581/DATA1_10  = p__arg0_0_8[10];
  assign \U581/DATA1_11  = p__arg0_0_8[11];
  assign \U580/DATA1_0  = p___constant_11x11xf32_0_8[0];
  assign \U580/DATA1_1  = p___constant_11x11xf32_0_8[1];
  assign \U580/DATA1_2  = p___constant_11x11xf32_0_8[2];
  assign \U580/DATA1_3  = p___constant_11x11xf32_0_8[3];
  assign \U580/DATA1_4  = p___constant_11x11xf32_0_8[4];
  assign \U580/DATA1_5  = p___constant_11x11xf32_0_8[5];
  assign \U580/DATA1_6  = p___constant_11x11xf32_0_8[6];
  assign \U580/DATA1_7  = p___constant_11x11xf32_0_8[7];
  assign \U580/DATA1_8  = p___constant_11x11xf32_0_8[8];
  assign \U580/DATA1_9  = p___constant_11x11xf32_0_8[9];
  assign \U580/DATA1_10  = p___constant_11x11xf32_0_8[10];
  assign \U580/DATA1_11  = p___constant_11x11xf32_0_8[11];
  assign \U576/DATA1_0  = p__arg0_0_9[0];
  assign \U576/DATA1_1  = p__arg0_0_9[1];
  assign \U576/DATA1_2  = p__arg0_0_9[2];
  assign \U576/DATA1_3  = p__arg0_0_9[3];
  assign \U576/DATA1_4  = p__arg0_0_9[4];
  assign \U576/DATA1_5  = p__arg0_0_9[5];
  assign \U576/DATA1_6  = p__arg0_0_9[6];
  assign \U576/DATA1_7  = p__arg0_0_9[7];
  assign \U576/DATA1_8  = p__arg0_0_9[8];
  assign \U576/DATA1_9  = p__arg0_0_9[9];
  assign \U576/DATA1_10  = p__arg0_0_9[10];
  assign \U576/DATA1_11  = p__arg0_0_9[11];
  assign \U575/DATA1_0  = p___constant_11x11xf32_0_9[0];
  assign \U575/DATA1_1  = p___constant_11x11xf32_0_9[1];
  assign \U575/DATA1_2  = p___constant_11x11xf32_0_9[2];
  assign \U575/DATA1_3  = p___constant_11x11xf32_0_9[3];
  assign \U575/DATA1_4  = p___constant_11x11xf32_0_9[4];
  assign \U575/DATA1_5  = p___constant_11x11xf32_0_9[5];
  assign \U575/DATA1_6  = p___constant_11x11xf32_0_9[6];
  assign \U575/DATA1_7  = p___constant_11x11xf32_0_9[7];
  assign \U575/DATA1_8  = p___constant_11x11xf32_0_9[8];
  assign \U575/DATA1_9  = p___constant_11x11xf32_0_9[9];
  assign \U575/DATA1_10  = p___constant_11x11xf32_0_9[10];
  assign \U575/DATA1_11  = p___constant_11x11xf32_0_9[11];
  assign \U571/DATA1_0  = p__arg0_0_10[0];
  assign \U571/DATA1_1  = p__arg0_0_10[1];
  assign \U571/DATA1_2  = p__arg0_0_10[2];
  assign \U571/DATA1_3  = p__arg0_0_10[3];
  assign \U571/DATA1_4  = p__arg0_0_10[4];
  assign \U571/DATA1_5  = p__arg0_0_10[5];
  assign \U571/DATA1_6  = p__arg0_0_10[6];
  assign \U571/DATA1_7  = p__arg0_0_10[7];
  assign \U571/DATA1_8  = p__arg0_0_10[8];
  assign \U571/DATA1_9  = p__arg0_0_10[9];
  assign \U571/DATA1_10  = p__arg0_0_10[10];
  assign \U571/DATA1_11  = p__arg0_0_10[11];
  assign \U570/DATA1_0  = p___constant_11x11xf32_0_10[0];
  assign \U570/DATA1_1  = p___constant_11x11xf32_0_10[1];
  assign \U570/DATA1_2  = p___constant_11x11xf32_0_10[2];
  assign \U570/DATA1_3  = p___constant_11x11xf32_0_10[3];
  assign \U570/DATA1_4  = p___constant_11x11xf32_0_10[4];
  assign \U570/DATA1_5  = p___constant_11x11xf32_0_10[5];
  assign \U570/DATA1_6  = p___constant_11x11xf32_0_10[6];
  assign \U570/DATA1_7  = p___constant_11x11xf32_0_10[7];
  assign \U570/DATA1_8  = p___constant_11x11xf32_0_10[8];
  assign \U570/DATA1_9  = p___constant_11x11xf32_0_10[9];
  assign \U570/DATA1_10  = p___constant_11x11xf32_0_10[10];
  assign \U570/DATA1_11  = p___constant_11x11xf32_0_10[11];
  assign \U565/DATA1_0  = p___constant_11xf32_0[0];
  assign \U565/DATA1_1  = p___constant_11xf32_0[1];
  assign \U565/DATA1_2  = p___constant_11xf32_0[2];
  assign \U565/DATA1_3  = p___constant_11xf32_0[3];
  assign \U565/DATA1_4  = p___constant_11xf32_0[4];
  assign \U565/DATA1_5  = p___constant_11xf32_0[5];
  assign \U565/DATA1_6  = p___constant_11xf32_0[6];
  assign \U565/DATA1_7  = p___constant_11xf32_0[7];
  assign \U565/DATA1_8  = p___constant_11xf32_0[8];
  assign \U565/DATA1_9  = p___constant_11xf32_0[9];
  assign \U565/DATA1_10  = p___constant_11xf32_0[10];
  assign \U565/DATA1_11  = p___constant_11xf32_0[11];
  assign \U553/DATA2_0  = p___constant_11x11xf32_1_0[0];
  assign \U553/DATA2_1  = p___constant_11x11xf32_1_0[1];
  assign \U553/DATA2_2  = p___constant_11x11xf32_1_0[2];
  assign \U553/DATA2_3  = p___constant_11x11xf32_1_0[3];
  assign \U553/DATA2_4  = p___constant_11x11xf32_1_0[4];
  assign \U553/DATA2_5  = p___constant_11x11xf32_1_0[5];
  assign \U553/DATA2_6  = p___constant_11x11xf32_1_0[6];
  assign \U553/DATA2_7  = p___constant_11x11xf32_1_0[7];
  assign \U553/DATA2_8  = p___constant_11x11xf32_1_0[8];
  assign \U553/DATA2_9  = p___constant_11x11xf32_1_0[9];
  assign \U553/DATA2_10  = p___constant_11x11xf32_1_0[10];
  assign \U553/DATA2_11  = p___constant_11x11xf32_1_0[11];
  assign \U553/DATA1_0  = p___constant_11x11xf32_1_1[0];
  assign \U553/DATA1_1  = p___constant_11x11xf32_1_1[1];
  assign \U553/DATA1_2  = p___constant_11x11xf32_1_1[2];
  assign \U553/DATA1_3  = p___constant_11x11xf32_1_1[3];
  assign \U553/DATA1_4  = p___constant_11x11xf32_1_1[4];
  assign \U553/DATA1_5  = p___constant_11x11xf32_1_1[5];
  assign \U553/DATA1_6  = p___constant_11x11xf32_1_1[6];
  assign \U553/DATA1_7  = p___constant_11x11xf32_1_1[7];
  assign \U553/DATA1_8  = p___constant_11x11xf32_1_1[8];
  assign \U553/DATA1_9  = p___constant_11x11xf32_1_1[9];
  assign \U553/DATA1_10  = p___constant_11x11xf32_1_1[10];
  assign \U553/DATA1_11  = p___constant_11x11xf32_1_1[11];
  assign \U548/DATA1_0  = p___constant_11x11xf32_1_2[0];
  assign \U548/DATA1_1  = p___constant_11x11xf32_1_2[1];
  assign \U548/DATA1_2  = p___constant_11x11xf32_1_2[2];
  assign \U548/DATA1_3  = p___constant_11x11xf32_1_2[3];
  assign \U548/DATA1_4  = p___constant_11x11xf32_1_2[4];
  assign \U548/DATA1_5  = p___constant_11x11xf32_1_2[5];
  assign \U548/DATA1_6  = p___constant_11x11xf32_1_2[6];
  assign \U548/DATA1_7  = p___constant_11x11xf32_1_2[7];
  assign \U548/DATA1_8  = p___constant_11x11xf32_1_2[8];
  assign \U548/DATA1_9  = p___constant_11x11xf32_1_2[9];
  assign \U548/DATA1_10  = p___constant_11x11xf32_1_2[10];
  assign \U548/DATA1_11  = p___constant_11x11xf32_1_2[11];
  assign \U543/DATA1_0  = p___constant_11x11xf32_1_3[0];
  assign \U543/DATA1_1  = p___constant_11x11xf32_1_3[1];
  assign \U543/DATA1_2  = p___constant_11x11xf32_1_3[2];
  assign \U543/DATA1_3  = p___constant_11x11xf32_1_3[3];
  assign \U543/DATA1_4  = p___constant_11x11xf32_1_3[4];
  assign \U543/DATA1_5  = p___constant_11x11xf32_1_3[5];
  assign \U543/DATA1_6  = p___constant_11x11xf32_1_3[6];
  assign \U543/DATA1_7  = p___constant_11x11xf32_1_3[7];
  assign \U543/DATA1_8  = p___constant_11x11xf32_1_3[8];
  assign \U543/DATA1_9  = p___constant_11x11xf32_1_3[9];
  assign \U543/DATA1_10  = p___constant_11x11xf32_1_3[10];
  assign \U543/DATA1_11  = p___constant_11x11xf32_1_3[11];
  assign \U538/DATA1_0  = p___constant_11x11xf32_1_4[0];
  assign \U538/DATA1_1  = p___constant_11x11xf32_1_4[1];
  assign \U538/DATA1_2  = p___constant_11x11xf32_1_4[2];
  assign \U538/DATA1_3  = p___constant_11x11xf32_1_4[3];
  assign \U538/DATA1_4  = p___constant_11x11xf32_1_4[4];
  assign \U538/DATA1_5  = p___constant_11x11xf32_1_4[5];
  assign \U538/DATA1_6  = p___constant_11x11xf32_1_4[6];
  assign \U538/DATA1_7  = p___constant_11x11xf32_1_4[7];
  assign \U538/DATA1_8  = p___constant_11x11xf32_1_4[8];
  assign \U538/DATA1_9  = p___constant_11x11xf32_1_4[9];
  assign \U538/DATA1_10  = p___constant_11x11xf32_1_4[10];
  assign \U538/DATA1_11  = p___constant_11x11xf32_1_4[11];
  assign \U533/DATA1_0  = p___constant_11x11xf32_1_5[0];
  assign \U533/DATA1_1  = p___constant_11x11xf32_1_5[1];
  assign \U533/DATA1_2  = p___constant_11x11xf32_1_5[2];
  assign \U533/DATA1_3  = p___constant_11x11xf32_1_5[3];
  assign \U533/DATA1_4  = p___constant_11x11xf32_1_5[4];
  assign \U533/DATA1_5  = p___constant_11x11xf32_1_5[5];
  assign \U533/DATA1_6  = p___constant_11x11xf32_1_5[6];
  assign \U533/DATA1_7  = p___constant_11x11xf32_1_5[7];
  assign \U533/DATA1_8  = p___constant_11x11xf32_1_5[8];
  assign \U533/DATA1_9  = p___constant_11x11xf32_1_5[9];
  assign \U533/DATA1_10  = p___constant_11x11xf32_1_5[10];
  assign \U533/DATA1_11  = p___constant_11x11xf32_1_5[11];
  assign \U528/DATA1_0  = p___constant_11x11xf32_1_6[0];
  assign \U528/DATA1_1  = p___constant_11x11xf32_1_6[1];
  assign \U528/DATA1_2  = p___constant_11x11xf32_1_6[2];
  assign \U528/DATA1_3  = p___constant_11x11xf32_1_6[3];
  assign \U528/DATA1_4  = p___constant_11x11xf32_1_6[4];
  assign \U528/DATA1_5  = p___constant_11x11xf32_1_6[5];
  assign \U528/DATA1_6  = p___constant_11x11xf32_1_6[6];
  assign \U528/DATA1_7  = p___constant_11x11xf32_1_6[7];
  assign \U528/DATA1_8  = p___constant_11x11xf32_1_6[8];
  assign \U528/DATA1_9  = p___constant_11x11xf32_1_6[9];
  assign \U528/DATA1_10  = p___constant_11x11xf32_1_6[10];
  assign \U528/DATA1_11  = p___constant_11x11xf32_1_6[11];
  assign \U523/DATA1_0  = p___constant_11x11xf32_1_7[0];
  assign \U523/DATA1_1  = p___constant_11x11xf32_1_7[1];
  assign \U523/DATA1_2  = p___constant_11x11xf32_1_7[2];
  assign \U523/DATA1_3  = p___constant_11x11xf32_1_7[3];
  assign \U523/DATA1_4  = p___constant_11x11xf32_1_7[4];
  assign \U523/DATA1_5  = p___constant_11x11xf32_1_7[5];
  assign \U523/DATA1_6  = p___constant_11x11xf32_1_7[6];
  assign \U523/DATA1_7  = p___constant_11x11xf32_1_7[7];
  assign \U523/DATA1_8  = p___constant_11x11xf32_1_7[8];
  assign \U523/DATA1_9  = p___constant_11x11xf32_1_7[9];
  assign \U523/DATA1_10  = p___constant_11x11xf32_1_7[10];
  assign \U523/DATA1_11  = p___constant_11x11xf32_1_7[11];
  assign \U518/DATA1_0  = p___constant_11x11xf32_1_8[0];
  assign \U518/DATA1_1  = p___constant_11x11xf32_1_8[1];
  assign \U518/DATA1_2  = p___constant_11x11xf32_1_8[2];
  assign \U518/DATA1_3  = p___constant_11x11xf32_1_8[3];
  assign \U518/DATA1_4  = p___constant_11x11xf32_1_8[4];
  assign \U518/DATA1_5  = p___constant_11x11xf32_1_8[5];
  assign \U518/DATA1_6  = p___constant_11x11xf32_1_8[6];
  assign \U518/DATA1_7  = p___constant_11x11xf32_1_8[7];
  assign \U518/DATA1_8  = p___constant_11x11xf32_1_8[8];
  assign \U518/DATA1_9  = p___constant_11x11xf32_1_8[9];
  assign \U518/DATA1_10  = p___constant_11x11xf32_1_8[10];
  assign \U518/DATA1_11  = p___constant_11x11xf32_1_8[11];
  assign \U513/DATA1_0  = p___constant_11x11xf32_1_9[0];
  assign \U513/DATA1_1  = p___constant_11x11xf32_1_9[1];
  assign \U513/DATA1_2  = p___constant_11x11xf32_1_9[2];
  assign \U513/DATA1_3  = p___constant_11x11xf32_1_9[3];
  assign \U513/DATA1_4  = p___constant_11x11xf32_1_9[4];
  assign \U513/DATA1_5  = p___constant_11x11xf32_1_9[5];
  assign \U513/DATA1_6  = p___constant_11x11xf32_1_9[6];
  assign \U513/DATA1_7  = p___constant_11x11xf32_1_9[7];
  assign \U513/DATA1_8  = p___constant_11x11xf32_1_9[8];
  assign \U513/DATA1_9  = p___constant_11x11xf32_1_9[9];
  assign \U513/DATA1_10  = p___constant_11x11xf32_1_9[10];
  assign \U513/DATA1_11  = p___constant_11x11xf32_1_9[11];
  assign \U508/DATA1_0  = p___constant_11x11xf32_1_10[0];
  assign \U508/DATA1_1  = p___constant_11x11xf32_1_10[1];
  assign \U508/DATA1_2  = p___constant_11x11xf32_1_10[2];
  assign \U508/DATA1_3  = p___constant_11x11xf32_1_10[3];
  assign \U508/DATA1_4  = p___constant_11x11xf32_1_10[4];
  assign \U508/DATA1_5  = p___constant_11x11xf32_1_10[5];
  assign \U508/DATA1_6  = p___constant_11x11xf32_1_10[6];
  assign \U508/DATA1_7  = p___constant_11x11xf32_1_10[7];
  assign \U508/DATA1_8  = p___constant_11x11xf32_1_10[8];
  assign \U508/DATA1_9  = p___constant_11x11xf32_1_10[9];
  assign \U508/DATA1_10  = p___constant_11x11xf32_1_10[10];
  assign \U508/DATA1_11  = p___constant_11x11xf32_1_10[11];
  assign \U503/DATA1_0  = p___constant_11xf32_1[0];
  assign \U503/DATA1_1  = p___constant_11xf32_1[1];
  assign \U503/DATA1_2  = p___constant_11xf32_1[2];
  assign \U503/DATA1_3  = p___constant_11xf32_1[3];
  assign \U503/DATA1_4  = p___constant_11xf32_1[4];
  assign \U503/DATA1_5  = p___constant_11xf32_1[5];
  assign \U503/DATA1_6  = p___constant_11xf32_1[6];
  assign \U503/DATA1_7  = p___constant_11xf32_1[7];
  assign \U503/DATA1_8  = p___constant_11xf32_1[8];
  assign \U503/DATA1_9  = p___constant_11xf32_1[9];
  assign \U503/DATA1_10  = p___constant_11xf32_1[10];
  assign \U503/DATA1_11  = p___constant_11xf32_1[11];
  assign \U500/DATA2_0  = p___constant_11x11xf32_2_0[0];
  assign \U500/DATA2_1  = p___constant_11x11xf32_2_0[1];
  assign \U500/DATA2_2  = p___constant_11x11xf32_2_0[2];
  assign \U500/DATA2_3  = p___constant_11x11xf32_2_0[3];
  assign \U500/DATA2_4  = p___constant_11x11xf32_2_0[4];
  assign \U500/DATA2_5  = p___constant_11x11xf32_2_0[5];
  assign \U500/DATA2_6  = p___constant_11x11xf32_2_0[6];
  assign \U500/DATA2_7  = p___constant_11x11xf32_2_0[7];
  assign \U500/DATA2_8  = p___constant_11x11xf32_2_0[8];
  assign \U500/DATA2_9  = p___constant_11x11xf32_2_0[9];
  assign \U500/DATA2_10  = p___constant_11x11xf32_2_0[10];
  assign \U500/DATA2_11  = p___constant_11x11xf32_2_0[11];
  assign \U500/DATA1_0  = p___constant_11x11xf32_2_1[0];
  assign \U500/DATA1_1  = p___constant_11x11xf32_2_1[1];
  assign \U500/DATA1_2  = p___constant_11x11xf32_2_1[2];
  assign \U500/DATA1_3  = p___constant_11x11xf32_2_1[3];
  assign \U500/DATA1_4  = p___constant_11x11xf32_2_1[4];
  assign \U500/DATA1_5  = p___constant_11x11xf32_2_1[5];
  assign \U500/DATA1_6  = p___constant_11x11xf32_2_1[6];
  assign \U500/DATA1_7  = p___constant_11x11xf32_2_1[7];
  assign \U500/DATA1_8  = p___constant_11x11xf32_2_1[8];
  assign \U500/DATA1_9  = p___constant_11x11xf32_2_1[9];
  assign \U500/DATA1_10  = p___constant_11x11xf32_2_1[10];
  assign \U500/DATA1_11  = p___constant_11x11xf32_2_1[11];
  assign \U495/DATA1_0  = p___constant_11x11xf32_2_2[0];
  assign \U495/DATA1_1  = p___constant_11x11xf32_2_2[1];
  assign \U495/DATA1_2  = p___constant_11x11xf32_2_2[2];
  assign \U495/DATA1_3  = p___constant_11x11xf32_2_2[3];
  assign \U495/DATA1_4  = p___constant_11x11xf32_2_2[4];
  assign \U495/DATA1_5  = p___constant_11x11xf32_2_2[5];
  assign \U495/DATA1_6  = p___constant_11x11xf32_2_2[6];
  assign \U495/DATA1_7  = p___constant_11x11xf32_2_2[7];
  assign \U495/DATA1_8  = p___constant_11x11xf32_2_2[8];
  assign \U495/DATA1_9  = p___constant_11x11xf32_2_2[9];
  assign \U495/DATA1_10  = p___constant_11x11xf32_2_2[10];
  assign \U495/DATA1_11  = p___constant_11x11xf32_2_2[11];
  assign \U490/DATA1_0  = p___constant_11x11xf32_2_3[0];
  assign \U490/DATA1_1  = p___constant_11x11xf32_2_3[1];
  assign \U490/DATA1_2  = p___constant_11x11xf32_2_3[2];
  assign \U490/DATA1_3  = p___constant_11x11xf32_2_3[3];
  assign \U490/DATA1_4  = p___constant_11x11xf32_2_3[4];
  assign \U490/DATA1_5  = p___constant_11x11xf32_2_3[5];
  assign \U490/DATA1_6  = p___constant_11x11xf32_2_3[6];
  assign \U490/DATA1_7  = p___constant_11x11xf32_2_3[7];
  assign \U490/DATA1_8  = p___constant_11x11xf32_2_3[8];
  assign \U490/DATA1_9  = p___constant_11x11xf32_2_3[9];
  assign \U490/DATA1_10  = p___constant_11x11xf32_2_3[10];
  assign \U490/DATA1_11  = p___constant_11x11xf32_2_3[11];
  assign \U485/DATA1_0  = p___constant_11x11xf32_2_4[0];
  assign \U485/DATA1_1  = p___constant_11x11xf32_2_4[1];
  assign \U485/DATA1_2  = p___constant_11x11xf32_2_4[2];
  assign \U485/DATA1_3  = p___constant_11x11xf32_2_4[3];
  assign \U485/DATA1_4  = p___constant_11x11xf32_2_4[4];
  assign \U485/DATA1_5  = p___constant_11x11xf32_2_4[5];
  assign \U485/DATA1_6  = p___constant_11x11xf32_2_4[6];
  assign \U485/DATA1_7  = p___constant_11x11xf32_2_4[7];
  assign \U485/DATA1_8  = p___constant_11x11xf32_2_4[8];
  assign \U485/DATA1_9  = p___constant_11x11xf32_2_4[9];
  assign \U485/DATA1_10  = p___constant_11x11xf32_2_4[10];
  assign \U485/DATA1_11  = p___constant_11x11xf32_2_4[11];
  assign \U480/DATA1_0  = p___constant_11x11xf32_2_5[0];
  assign \U480/DATA1_1  = p___constant_11x11xf32_2_5[1];
  assign \U480/DATA1_2  = p___constant_11x11xf32_2_5[2];
  assign \U480/DATA1_3  = p___constant_11x11xf32_2_5[3];
  assign \U480/DATA1_4  = p___constant_11x11xf32_2_5[4];
  assign \U480/DATA1_5  = p___constant_11x11xf32_2_5[5];
  assign \U480/DATA1_6  = p___constant_11x11xf32_2_5[6];
  assign \U480/DATA1_7  = p___constant_11x11xf32_2_5[7];
  assign \U480/DATA1_8  = p___constant_11x11xf32_2_5[8];
  assign \U480/DATA1_9  = p___constant_11x11xf32_2_5[9];
  assign \U480/DATA1_10  = p___constant_11x11xf32_2_5[10];
  assign \U480/DATA1_11  = p___constant_11x11xf32_2_5[11];
  assign \U475/DATA1_0  = p___constant_11x11xf32_2_6[0];
  assign \U475/DATA1_1  = p___constant_11x11xf32_2_6[1];
  assign \U475/DATA1_2  = p___constant_11x11xf32_2_6[2];
  assign \U475/DATA1_3  = p___constant_11x11xf32_2_6[3];
  assign \U475/DATA1_4  = p___constant_11x11xf32_2_6[4];
  assign \U475/DATA1_5  = p___constant_11x11xf32_2_6[5];
  assign \U475/DATA1_6  = p___constant_11x11xf32_2_6[6];
  assign \U475/DATA1_7  = p___constant_11x11xf32_2_6[7];
  assign \U475/DATA1_8  = p___constant_11x11xf32_2_6[8];
  assign \U475/DATA1_9  = p___constant_11x11xf32_2_6[9];
  assign \U475/DATA1_10  = p___constant_11x11xf32_2_6[10];
  assign \U475/DATA1_11  = p___constant_11x11xf32_2_6[11];
  assign \U470/DATA1_0  = p___constant_11x11xf32_2_7[0];
  assign \U470/DATA1_1  = p___constant_11x11xf32_2_7[1];
  assign \U470/DATA1_2  = p___constant_11x11xf32_2_7[2];
  assign \U470/DATA1_3  = p___constant_11x11xf32_2_7[3];
  assign \U470/DATA1_4  = p___constant_11x11xf32_2_7[4];
  assign \U470/DATA1_5  = p___constant_11x11xf32_2_7[5];
  assign \U470/DATA1_6  = p___constant_11x11xf32_2_7[6];
  assign \U470/DATA1_7  = p___constant_11x11xf32_2_7[7];
  assign \U470/DATA1_8  = p___constant_11x11xf32_2_7[8];
  assign \U470/DATA1_9  = p___constant_11x11xf32_2_7[9];
  assign \U470/DATA1_10  = p___constant_11x11xf32_2_7[10];
  assign \U470/DATA1_11  = p___constant_11x11xf32_2_7[11];
  assign \U465/DATA1_0  = p___constant_11x11xf32_2_8[0];
  assign \U465/DATA1_1  = p___constant_11x11xf32_2_8[1];
  assign \U465/DATA1_2  = p___constant_11x11xf32_2_8[2];
  assign \U465/DATA1_3  = p___constant_11x11xf32_2_8[3];
  assign \U465/DATA1_4  = p___constant_11x11xf32_2_8[4];
  assign \U465/DATA1_5  = p___constant_11x11xf32_2_8[5];
  assign \U465/DATA1_6  = p___constant_11x11xf32_2_8[6];
  assign \U465/DATA1_7  = p___constant_11x11xf32_2_8[7];
  assign \U465/DATA1_8  = p___constant_11x11xf32_2_8[8];
  assign \U465/DATA1_9  = p___constant_11x11xf32_2_8[9];
  assign \U465/DATA1_10  = p___constant_11x11xf32_2_8[10];
  assign \U465/DATA1_11  = p___constant_11x11xf32_2_8[11];
  assign \U460/DATA1_0  = p___constant_11x11xf32_2_9[0];
  assign \U460/DATA1_1  = p___constant_11x11xf32_2_9[1];
  assign \U460/DATA1_2  = p___constant_11x11xf32_2_9[2];
  assign \U460/DATA1_3  = p___constant_11x11xf32_2_9[3];
  assign \U460/DATA1_4  = p___constant_11x11xf32_2_9[4];
  assign \U460/DATA1_5  = p___constant_11x11xf32_2_9[5];
  assign \U460/DATA1_6  = p___constant_11x11xf32_2_9[6];
  assign \U460/DATA1_7  = p___constant_11x11xf32_2_9[7];
  assign \U460/DATA1_8  = p___constant_11x11xf32_2_9[8];
  assign \U460/DATA1_9  = p___constant_11x11xf32_2_9[9];
  assign \U460/DATA1_10  = p___constant_11x11xf32_2_9[10];
  assign \U460/DATA1_11  = p___constant_11x11xf32_2_9[11];
  assign \U455/DATA1_0  = p___constant_11x11xf32_2_10[0];
  assign \U455/DATA1_1  = p___constant_11x11xf32_2_10[1];
  assign \U455/DATA1_2  = p___constant_11x11xf32_2_10[2];
  assign \U455/DATA1_3  = p___constant_11x11xf32_2_10[3];
  assign \U455/DATA1_4  = p___constant_11x11xf32_2_10[4];
  assign \U455/DATA1_5  = p___constant_11x11xf32_2_10[5];
  assign \U455/DATA1_6  = p___constant_11x11xf32_2_10[6];
  assign \U455/DATA1_7  = p___constant_11x11xf32_2_10[7];
  assign \U455/DATA1_8  = p___constant_11x11xf32_2_10[8];
  assign \U455/DATA1_9  = p___constant_11x11xf32_2_10[9];
  assign \U455/DATA1_10  = p___constant_11x11xf32_2_10[10];
  assign \U455/DATA1_11  = p___constant_11x11xf32_2_10[11];
  assign \U450/DATA1_0  = p___constant_11xf32_2[0];
  assign \U450/DATA1_1  = p___constant_11xf32_2[1];
  assign \U450/DATA1_2  = p___constant_11xf32_2[2];
  assign \U450/DATA1_3  = p___constant_11xf32_2[3];
  assign \U450/DATA1_4  = p___constant_11xf32_2[4];
  assign \U450/DATA1_5  = p___constant_11xf32_2[5];
  assign \U450/DATA1_6  = p___constant_11xf32_2[6];
  assign \U450/DATA1_7  = p___constant_11xf32_2[7];
  assign \U450/DATA1_8  = p___constant_11xf32_2[8];
  assign \U450/DATA1_9  = p___constant_11xf32_2[9];
  assign \U450/DATA1_10  = p___constant_11xf32_2[10];
  assign \U450/DATA1_11  = p___constant_11xf32_2[11];
  assign \U444/DATA2_0  = p___constant_11x11xf32_3_0[0];
  assign \U444/DATA2_1  = p___constant_11x11xf32_3_0[1];
  assign \U444/DATA2_2  = p___constant_11x11xf32_3_0[2];
  assign \U444/DATA2_3  = p___constant_11x11xf32_3_0[3];
  assign \U444/DATA2_4  = p___constant_11x11xf32_3_0[4];
  assign \U444/DATA2_5  = p___constant_11x11xf32_3_0[5];
  assign \U444/DATA2_6  = p___constant_11x11xf32_3_0[6];
  assign \U444/DATA2_7  = p___constant_11x11xf32_3_0[7];
  assign \U444/DATA2_8  = p___constant_11x11xf32_3_0[8];
  assign \U444/DATA2_9  = p___constant_11x11xf32_3_0[9];
  assign \U444/DATA2_10  = p___constant_11x11xf32_3_0[10];
  assign \U444/DATA2_11  = p___constant_11x11xf32_3_0[11];
  assign \U444/DATA1_0  = p___constant_11x11xf32_3_1[0];
  assign \U444/DATA1_1  = p___constant_11x11xf32_3_1[1];
  assign \U444/DATA1_2  = p___constant_11x11xf32_3_1[2];
  assign \U444/DATA1_3  = p___constant_11x11xf32_3_1[3];
  assign \U444/DATA1_4  = p___constant_11x11xf32_3_1[4];
  assign \U444/DATA1_5  = p___constant_11x11xf32_3_1[5];
  assign \U444/DATA1_6  = p___constant_11x11xf32_3_1[6];
  assign \U444/DATA1_7  = p___constant_11x11xf32_3_1[7];
  assign \U444/DATA1_8  = p___constant_11x11xf32_3_1[8];
  assign \U444/DATA1_9  = p___constant_11x11xf32_3_1[9];
  assign \U444/DATA1_10  = p___constant_11x11xf32_3_1[10];
  assign \U444/DATA1_11  = p___constant_11x11xf32_3_1[11];
  assign \U439/DATA1_0  = p___constant_11x11xf32_3_2[0];
  assign \U439/DATA1_1  = p___constant_11x11xf32_3_2[1];
  assign \U439/DATA1_2  = p___constant_11x11xf32_3_2[2];
  assign \U439/DATA1_3  = p___constant_11x11xf32_3_2[3];
  assign \U439/DATA1_4  = p___constant_11x11xf32_3_2[4];
  assign \U439/DATA1_5  = p___constant_11x11xf32_3_2[5];
  assign \U439/DATA1_6  = p___constant_11x11xf32_3_2[6];
  assign \U439/DATA1_7  = p___constant_11x11xf32_3_2[7];
  assign \U439/DATA1_8  = p___constant_11x11xf32_3_2[8];
  assign \U439/DATA1_9  = p___constant_11x11xf32_3_2[9];
  assign \U439/DATA1_10  = p___constant_11x11xf32_3_2[10];
  assign \U439/DATA1_11  = p___constant_11x11xf32_3_2[11];
  assign \U434/DATA1_0  = p___constant_11x11xf32_3_3[0];
  assign \U434/DATA1_1  = p___constant_11x11xf32_3_3[1];
  assign \U434/DATA1_2  = p___constant_11x11xf32_3_3[2];
  assign \U434/DATA1_3  = p___constant_11x11xf32_3_3[3];
  assign \U434/DATA1_4  = p___constant_11x11xf32_3_3[4];
  assign \U434/DATA1_5  = p___constant_11x11xf32_3_3[5];
  assign \U434/DATA1_6  = p___constant_11x11xf32_3_3[6];
  assign \U434/DATA1_7  = p___constant_11x11xf32_3_3[7];
  assign \U434/DATA1_8  = p___constant_11x11xf32_3_3[8];
  assign \U434/DATA1_9  = p___constant_11x11xf32_3_3[9];
  assign \U434/DATA1_10  = p___constant_11x11xf32_3_3[10];
  assign \U434/DATA1_11  = p___constant_11x11xf32_3_3[11];
  assign \U429/DATA1_0  = p___constant_11x11xf32_3_4[0];
  assign \U429/DATA1_1  = p___constant_11x11xf32_3_4[1];
  assign \U429/DATA1_2  = p___constant_11x11xf32_3_4[2];
  assign \U429/DATA1_3  = p___constant_11x11xf32_3_4[3];
  assign \U429/DATA1_4  = p___constant_11x11xf32_3_4[4];
  assign \U429/DATA1_5  = p___constant_11x11xf32_3_4[5];
  assign \U429/DATA1_6  = p___constant_11x11xf32_3_4[6];
  assign \U429/DATA1_7  = p___constant_11x11xf32_3_4[7];
  assign \U429/DATA1_8  = p___constant_11x11xf32_3_4[8];
  assign \U429/DATA1_9  = p___constant_11x11xf32_3_4[9];
  assign \U429/DATA1_10  = p___constant_11x11xf32_3_4[10];
  assign \U429/DATA1_11  = p___constant_11x11xf32_3_4[11];
  assign \U424/DATA1_0  = p___constant_11x11xf32_3_5[0];
  assign \U424/DATA1_1  = p___constant_11x11xf32_3_5[1];
  assign \U424/DATA1_2  = p___constant_11x11xf32_3_5[2];
  assign \U424/DATA1_3  = p___constant_11x11xf32_3_5[3];
  assign \U424/DATA1_4  = p___constant_11x11xf32_3_5[4];
  assign \U424/DATA1_5  = p___constant_11x11xf32_3_5[5];
  assign \U424/DATA1_6  = p___constant_11x11xf32_3_5[6];
  assign \U424/DATA1_7  = p___constant_11x11xf32_3_5[7];
  assign \U424/DATA1_8  = p___constant_11x11xf32_3_5[8];
  assign \U424/DATA1_9  = p___constant_11x11xf32_3_5[9];
  assign \U424/DATA1_10  = p___constant_11x11xf32_3_5[10];
  assign \U424/DATA1_11  = p___constant_11x11xf32_3_5[11];
  assign \U419/DATA1_0  = p___constant_11x11xf32_3_6[0];
  assign \U419/DATA1_1  = p___constant_11x11xf32_3_6[1];
  assign \U419/DATA1_2  = p___constant_11x11xf32_3_6[2];
  assign \U419/DATA1_3  = p___constant_11x11xf32_3_6[3];
  assign \U419/DATA1_4  = p___constant_11x11xf32_3_6[4];
  assign \U419/DATA1_5  = p___constant_11x11xf32_3_6[5];
  assign \U419/DATA1_6  = p___constant_11x11xf32_3_6[6];
  assign \U419/DATA1_7  = p___constant_11x11xf32_3_6[7];
  assign \U419/DATA1_8  = p___constant_11x11xf32_3_6[8];
  assign \U419/DATA1_9  = p___constant_11x11xf32_3_6[9];
  assign \U419/DATA1_10  = p___constant_11x11xf32_3_6[10];
  assign \U419/DATA1_11  = p___constant_11x11xf32_3_6[11];
  assign \U414/DATA1_0  = p___constant_11x11xf32_3_7[0];
  assign \U414/DATA1_1  = p___constant_11x11xf32_3_7[1];
  assign \U414/DATA1_2  = p___constant_11x11xf32_3_7[2];
  assign \U414/DATA1_3  = p___constant_11x11xf32_3_7[3];
  assign \U414/DATA1_4  = p___constant_11x11xf32_3_7[4];
  assign \U414/DATA1_5  = p___constant_11x11xf32_3_7[5];
  assign \U414/DATA1_6  = p___constant_11x11xf32_3_7[6];
  assign \U414/DATA1_7  = p___constant_11x11xf32_3_7[7];
  assign \U414/DATA1_8  = p___constant_11x11xf32_3_7[8];
  assign \U414/DATA1_9  = p___constant_11x11xf32_3_7[9];
  assign \U414/DATA1_10  = p___constant_11x11xf32_3_7[10];
  assign \U414/DATA1_11  = p___constant_11x11xf32_3_7[11];
  assign \U409/DATA1_0  = p___constant_11x11xf32_3_8[0];
  assign \U409/DATA1_1  = p___constant_11x11xf32_3_8[1];
  assign \U409/DATA1_2  = p___constant_11x11xf32_3_8[2];
  assign \U409/DATA1_3  = p___constant_11x11xf32_3_8[3];
  assign \U409/DATA1_4  = p___constant_11x11xf32_3_8[4];
  assign \U409/DATA1_5  = p___constant_11x11xf32_3_8[5];
  assign \U409/DATA1_6  = p___constant_11x11xf32_3_8[6];
  assign \U409/DATA1_7  = p___constant_11x11xf32_3_8[7];
  assign \U409/DATA1_8  = p___constant_11x11xf32_3_8[8];
  assign \U409/DATA1_9  = p___constant_11x11xf32_3_8[9];
  assign \U409/DATA1_10  = p___constant_11x11xf32_3_8[10];
  assign \U409/DATA1_11  = p___constant_11x11xf32_3_8[11];
  assign \U404/DATA1_0  = p___constant_11x11xf32_3_9[0];
  assign \U404/DATA1_1  = p___constant_11x11xf32_3_9[1];
  assign \U404/DATA1_2  = p___constant_11x11xf32_3_9[2];
  assign \U404/DATA1_3  = p___constant_11x11xf32_3_9[3];
  assign \U404/DATA1_4  = p___constant_11x11xf32_3_9[4];
  assign \U404/DATA1_5  = p___constant_11x11xf32_3_9[5];
  assign \U404/DATA1_6  = p___constant_11x11xf32_3_9[6];
  assign \U404/DATA1_7  = p___constant_11x11xf32_3_9[7];
  assign \U404/DATA1_8  = p___constant_11x11xf32_3_9[8];
  assign \U404/DATA1_9  = p___constant_11x11xf32_3_9[9];
  assign \U404/DATA1_10  = p___constant_11x11xf32_3_9[10];
  assign \U404/DATA1_11  = p___constant_11x11xf32_3_9[11];
  assign \U399/DATA1_0  = p___constant_11x11xf32_3_10[0];
  assign \U399/DATA1_1  = p___constant_11x11xf32_3_10[1];
  assign \U399/DATA1_2  = p___constant_11x11xf32_3_10[2];
  assign \U399/DATA1_3  = p___constant_11x11xf32_3_10[3];
  assign \U399/DATA1_4  = p___constant_11x11xf32_3_10[4];
  assign \U399/DATA1_5  = p___constant_11x11xf32_3_10[5];
  assign \U399/DATA1_6  = p___constant_11x11xf32_3_10[6];
  assign \U399/DATA1_7  = p___constant_11x11xf32_3_10[7];
  assign \U399/DATA1_8  = p___constant_11x11xf32_3_10[8];
  assign \U399/DATA1_9  = p___constant_11x11xf32_3_10[9];
  assign \U399/DATA1_10  = p___constant_11x11xf32_3_10[10];
  assign \U399/DATA1_11  = p___constant_11x11xf32_3_10[11];
  assign \U394/DATA1_0  = p___constant_11xf32_3[0];
  assign \U394/DATA1_1  = p___constant_11xf32_3[1];
  assign \U394/DATA1_2  = p___constant_11xf32_3[2];
  assign \U394/DATA1_3  = p___constant_11xf32_3[3];
  assign \U394/DATA1_4  = p___constant_11xf32_3[4];
  assign \U394/DATA1_5  = p___constant_11xf32_3[5];
  assign \U394/DATA1_6  = p___constant_11xf32_3[6];
  assign \U394/DATA1_7  = p___constant_11xf32_3[7];
  assign \U394/DATA1_8  = p___constant_11xf32_3[8];
  assign \U394/DATA1_9  = p___constant_11xf32_3[9];
  assign \U394/DATA1_10  = p___constant_11xf32_3[10];
  assign \U394/DATA1_11  = p___constant_11xf32_3[11];
  assign \U391/DATA2_0  = p___constant_11x11xf32_4_0[0];
  assign \U391/DATA2_1  = p___constant_11x11xf32_4_0[1];
  assign \U391/DATA2_2  = p___constant_11x11xf32_4_0[2];
  assign \U391/DATA2_3  = p___constant_11x11xf32_4_0[3];
  assign \U391/DATA2_4  = p___constant_11x11xf32_4_0[4];
  assign \U391/DATA2_5  = p___constant_11x11xf32_4_0[5];
  assign \U391/DATA2_6  = p___constant_11x11xf32_4_0[6];
  assign \U391/DATA2_7  = p___constant_11x11xf32_4_0[7];
  assign \U391/DATA2_8  = p___constant_11x11xf32_4_0[8];
  assign \U391/DATA2_9  = p___constant_11x11xf32_4_0[9];
  assign \U391/DATA2_10  = p___constant_11x11xf32_4_0[10];
  assign \U391/DATA2_11  = p___constant_11x11xf32_4_0[11];
  assign \U391/DATA1_0  = p___constant_11x11xf32_4_1[0];
  assign \U391/DATA1_1  = p___constant_11x11xf32_4_1[1];
  assign \U391/DATA1_2  = p___constant_11x11xf32_4_1[2];
  assign \U391/DATA1_3  = p___constant_11x11xf32_4_1[3];
  assign \U391/DATA1_4  = p___constant_11x11xf32_4_1[4];
  assign \U391/DATA1_5  = p___constant_11x11xf32_4_1[5];
  assign \U391/DATA1_6  = p___constant_11x11xf32_4_1[6];
  assign \U391/DATA1_7  = p___constant_11x11xf32_4_1[7];
  assign \U391/DATA1_8  = p___constant_11x11xf32_4_1[8];
  assign \U391/DATA1_9  = p___constant_11x11xf32_4_1[9];
  assign \U391/DATA1_10  = p___constant_11x11xf32_4_1[10];
  assign \U391/DATA1_11  = p___constant_11x11xf32_4_1[11];
  assign \U386/DATA1_0  = p___constant_11x11xf32_4_2[0];
  assign \U386/DATA1_1  = p___constant_11x11xf32_4_2[1];
  assign \U386/DATA1_2  = p___constant_11x11xf32_4_2[2];
  assign \U386/DATA1_3  = p___constant_11x11xf32_4_2[3];
  assign \U386/DATA1_4  = p___constant_11x11xf32_4_2[4];
  assign \U386/DATA1_5  = p___constant_11x11xf32_4_2[5];
  assign \U386/DATA1_6  = p___constant_11x11xf32_4_2[6];
  assign \U386/DATA1_7  = p___constant_11x11xf32_4_2[7];
  assign \U386/DATA1_8  = p___constant_11x11xf32_4_2[8];
  assign \U386/DATA1_9  = p___constant_11x11xf32_4_2[9];
  assign \U386/DATA1_10  = p___constant_11x11xf32_4_2[10];
  assign \U386/DATA1_11  = p___constant_11x11xf32_4_2[11];
  assign \U381/DATA1_0  = p___constant_11x11xf32_4_3[0];
  assign \U381/DATA1_1  = p___constant_11x11xf32_4_3[1];
  assign \U381/DATA1_2  = p___constant_11x11xf32_4_3[2];
  assign \U381/DATA1_3  = p___constant_11x11xf32_4_3[3];
  assign \U381/DATA1_4  = p___constant_11x11xf32_4_3[4];
  assign \U381/DATA1_5  = p___constant_11x11xf32_4_3[5];
  assign \U381/DATA1_6  = p___constant_11x11xf32_4_3[6];
  assign \U381/DATA1_7  = p___constant_11x11xf32_4_3[7];
  assign \U381/DATA1_8  = p___constant_11x11xf32_4_3[8];
  assign \U381/DATA1_9  = p___constant_11x11xf32_4_3[9];
  assign \U381/DATA1_10  = p___constant_11x11xf32_4_3[10];
  assign \U381/DATA1_11  = p___constant_11x11xf32_4_3[11];
  assign \U376/DATA1_0  = p___constant_11x11xf32_4_4[0];
  assign \U376/DATA1_1  = p___constant_11x11xf32_4_4[1];
  assign \U376/DATA1_2  = p___constant_11x11xf32_4_4[2];
  assign \U376/DATA1_3  = p___constant_11x11xf32_4_4[3];
  assign \U376/DATA1_4  = p___constant_11x11xf32_4_4[4];
  assign \U376/DATA1_5  = p___constant_11x11xf32_4_4[5];
  assign \U376/DATA1_6  = p___constant_11x11xf32_4_4[6];
  assign \U376/DATA1_7  = p___constant_11x11xf32_4_4[7];
  assign \U376/DATA1_8  = p___constant_11x11xf32_4_4[8];
  assign \U376/DATA1_9  = p___constant_11x11xf32_4_4[9];
  assign \U376/DATA1_10  = p___constant_11x11xf32_4_4[10];
  assign \U376/DATA1_11  = p___constant_11x11xf32_4_4[11];
  assign \U371/DATA1_0  = p___constant_11x11xf32_4_5[0];
  assign \U371/DATA1_1  = p___constant_11x11xf32_4_5[1];
  assign \U371/DATA1_2  = p___constant_11x11xf32_4_5[2];
  assign \U371/DATA1_3  = p___constant_11x11xf32_4_5[3];
  assign \U371/DATA1_4  = p___constant_11x11xf32_4_5[4];
  assign \U371/DATA1_5  = p___constant_11x11xf32_4_5[5];
  assign \U371/DATA1_6  = p___constant_11x11xf32_4_5[6];
  assign \U371/DATA1_7  = p___constant_11x11xf32_4_5[7];
  assign \U371/DATA1_8  = p___constant_11x11xf32_4_5[8];
  assign \U371/DATA1_9  = p___constant_11x11xf32_4_5[9];
  assign \U371/DATA1_10  = p___constant_11x11xf32_4_5[10];
  assign \U371/DATA1_11  = p___constant_11x11xf32_4_5[11];
  assign \U366/DATA1_0  = p___constant_11x11xf32_4_6[0];
  assign \U366/DATA1_1  = p___constant_11x11xf32_4_6[1];
  assign \U366/DATA1_2  = p___constant_11x11xf32_4_6[2];
  assign \U366/DATA1_3  = p___constant_11x11xf32_4_6[3];
  assign \U366/DATA1_4  = p___constant_11x11xf32_4_6[4];
  assign \U366/DATA1_5  = p___constant_11x11xf32_4_6[5];
  assign \U366/DATA1_6  = p___constant_11x11xf32_4_6[6];
  assign \U366/DATA1_7  = p___constant_11x11xf32_4_6[7];
  assign \U366/DATA1_8  = p___constant_11x11xf32_4_6[8];
  assign \U366/DATA1_9  = p___constant_11x11xf32_4_6[9];
  assign \U366/DATA1_10  = p___constant_11x11xf32_4_6[10];
  assign \U366/DATA1_11  = p___constant_11x11xf32_4_6[11];
  assign \U361/DATA1_3  = p___constant_11x11xf32_4_7[3];
  assign \U361/DATA1_4  = p___constant_11x11xf32_4_7[4];
  assign \U361/DATA1_5  = p___constant_11x11xf32_4_7[5];
  assign \U361/DATA1_6  = p___constant_11x11xf32_4_7[6];
  assign \U361/DATA1_7  = p___constant_11x11xf32_4_7[7];
  assign \U361/DATA1_8  = p___constant_11x11xf32_4_7[8];
  assign \U361/DATA1_9  = p___constant_11x11xf32_4_7[9];
  assign \U361/DATA1_10  = p___constant_11x11xf32_4_7[10];
  assign \U361/DATA1_11  = p___constant_11x11xf32_4_7[11];
  assign \U356/DATA1_1  = p___constant_11x11xf32_4_8[1];
  assign \U356/DATA1_2  = p___constant_11x11xf32_4_8[2];
  assign \U356/DATA1_3  = p___constant_11x11xf32_4_8[3];
  assign \U356/DATA1_4  = p___constant_11x11xf32_4_8[4];
  assign \U356/DATA1_5  = p___constant_11x11xf32_4_8[5];
  assign \U356/DATA1_6  = p___constant_11x11xf32_4_8[6];
  assign \U356/DATA1_7  = p___constant_11x11xf32_4_8[7];
  assign \U356/DATA1_8  = p___constant_11x11xf32_4_8[8];
  assign \U356/DATA1_9  = p___constant_11x11xf32_4_8[9];
  assign \U356/DATA1_10  = p___constant_11x11xf32_4_8[10];
  assign \U356/DATA1_11  = p___constant_11x11xf32_4_8[11];
  assign \U351/DATA1_1  = p___constant_11x11xf32_4_9[1];
  assign \U351/DATA1_2  = p___constant_11x11xf32_4_9[2];
  assign \U351/DATA1_3  = p___constant_11x11xf32_4_9[3];
  assign \U351/DATA1_4  = p___constant_11x11xf32_4_9[4];
  assign \U351/DATA1_5  = p___constant_11x11xf32_4_9[5];
  assign \U351/DATA1_6  = p___constant_11x11xf32_4_9[6];
  assign \U351/DATA1_7  = p___constant_11x11xf32_4_9[7];
  assign \U351/DATA1_8  = p___constant_11x11xf32_4_9[8];
  assign \U351/DATA1_9  = p___constant_11x11xf32_4_9[9];
  assign \U351/DATA1_10  = p___constant_11x11xf32_4_9[10];
  assign \U351/DATA1_11  = p___constant_11x11xf32_4_9[11];
  assign \U346/DATA1_5  = p___constant_11x11xf32_4_10[5];
  assign \U346/DATA1_6  = p___constant_11x11xf32_4_10[6];
  assign \U346/DATA1_7  = p___constant_11x11xf32_4_10[7];
  assign \U346/DATA1_8  = p___constant_11x11xf32_4_10[8];
  assign \U346/DATA1_9  = p___constant_11x11xf32_4_10[9];
  assign \U346/DATA1_10  = p___constant_11x11xf32_4_10[10];
  assign \U346/DATA1_11  = p___constant_11x11xf32_4_10[11];
  assign \U341/DATA1_1  = p___constant_11xf32_4[1];
  assign \U341/DATA1_2  = p___constant_11xf32_4[2];
  assign \U341/DATA1_3  = p___constant_11xf32_4[3];
  assign \U341/DATA1_4  = p___constant_11xf32_4[4];
  assign \U341/DATA1_5  = p___constant_11xf32_4[5];
  assign \U341/DATA1_6  = p___constant_11xf32_4[6];
  assign \U341/DATA1_7  = p___constant_11xf32_4[7];
  assign \U341/DATA1_8  = p___constant_11xf32_4[8];
  assign \U341/DATA1_9  = p___constant_11xf32_4[9];
  assign \U341/DATA1_10  = p___constant_11xf32_4[10];
  assign \U341/DATA1_11  = p___constant_11xf32_4[11];
  assign \U332/DATA2_1  = p___constant_11x11xf32_5_0[1];
  assign \U332/DATA2_2  = p___constant_11x11xf32_5_0[2];
  assign \U332/DATA2_3  = p___constant_11x11xf32_5_0[3];
  assign \U332/DATA2_4  = p___constant_11x11xf32_5_0[4];
  assign \U332/DATA2_5  = p___constant_11x11xf32_5_0[5];
  assign \U332/DATA2_6  = p___constant_11x11xf32_5_0[6];
  assign \U332/DATA2_7  = p___constant_11x11xf32_5_0[7];
  assign \U332/DATA2_8  = p___constant_11x11xf32_5_0[8];
  assign \U332/DATA2_9  = p___constant_11x11xf32_5_0[9];
  assign \U332/DATA2_10  = p___constant_11x11xf32_5_0[10];
  assign \U332/DATA2_11  = p___constant_11x11xf32_5_0[11];
  assign \U332/DATA1_1  = p___constant_11x11xf32_5_1[1];
  assign \U332/DATA1_2  = p___constant_11x11xf32_5_1[2];
  assign \U332/DATA1_3  = p___constant_11x11xf32_5_1[3];
  assign \U332/DATA1_4  = p___constant_11x11xf32_5_1[4];
  assign \U332/DATA1_5  = p___constant_11x11xf32_5_1[5];
  assign \U332/DATA1_6  = p___constant_11x11xf32_5_1[6];
  assign \U332/DATA1_7  = p___constant_11x11xf32_5_1[7];
  assign \U332/DATA1_8  = p___constant_11x11xf32_5_1[8];
  assign \U332/DATA1_9  = p___constant_11x11xf32_5_1[9];
  assign \U332/DATA1_10  = p___constant_11x11xf32_5_1[10];
  assign \U332/DATA1_11  = p___constant_11x11xf32_5_1[11];
  assign \U327/DATA1_2  = p___constant_11x11xf32_5_2[2];
  assign \U327/DATA1_3  = p___constant_11x11xf32_5_2[3];
  assign \U327/DATA1_4  = p___constant_11x11xf32_5_2[4];
  assign \U327/DATA1_5  = p___constant_11x11xf32_5_2[5];
  assign \U327/DATA1_6  = p___constant_11x11xf32_5_2[6];
  assign \U327/DATA1_7  = p___constant_11x11xf32_5_2[7];
  assign \U327/DATA1_8  = p___constant_11x11xf32_5_2[8];
  assign \U327/DATA1_9  = p___constant_11x11xf32_5_2[9];
  assign \U327/DATA1_10  = p___constant_11x11xf32_5_2[10];
  assign \U327/DATA1_11  = p___constant_11x11xf32_5_2[11];
  assign \U322/DATA1_3  = p___constant_11x11xf32_5_3[3];
  assign \U322/DATA1_4  = p___constant_11x11xf32_5_3[4];
  assign \U322/DATA1_5  = p___constant_11x11xf32_5_3[5];
  assign \U322/DATA1_6  = p___constant_11x11xf32_5_3[6];
  assign \U322/DATA1_7  = p___constant_11x11xf32_5_3[7];
  assign \U322/DATA1_8  = p___constant_11x11xf32_5_3[8];
  assign \U322/DATA1_9  = p___constant_11x11xf32_5_3[9];
  assign \U322/DATA1_10  = p___constant_11x11xf32_5_3[10];
  assign \U322/DATA1_11  = p___constant_11x11xf32_5_3[11];
  assign \U317/DATA1_1  = p___constant_11x11xf32_5_4[1];
  assign \U317/DATA1_2  = p___constant_11x11xf32_5_4[2];
  assign \U317/DATA1_3  = p___constant_11x11xf32_5_4[3];
  assign \U317/DATA1_4  = p___constant_11x11xf32_5_4[4];
  assign \U317/DATA1_5  = p___constant_11x11xf32_5_4[5];
  assign \U317/DATA1_6  = p___constant_11x11xf32_5_4[6];
  assign \U317/DATA1_7  = p___constant_11x11xf32_5_4[7];
  assign \U317/DATA1_8  = p___constant_11x11xf32_5_4[8];
  assign \U317/DATA1_9  = p___constant_11x11xf32_5_4[9];
  assign \U317/DATA1_10  = p___constant_11x11xf32_5_4[10];
  assign \U317/DATA1_11  = p___constant_11x11xf32_5_4[11];
  assign \U312/DATA1_1  = p___constant_11x11xf32_5_5[1];
  assign \U312/DATA1_2  = p___constant_11x11xf32_5_5[2];
  assign \U312/DATA1_3  = p___constant_11x11xf32_5_5[3];
  assign \U312/DATA1_4  = p___constant_11x11xf32_5_5[4];
  assign \U312/DATA1_5  = p___constant_11x11xf32_5_5[5];
  assign \U312/DATA1_6  = p___constant_11x11xf32_5_5[6];
  assign \U312/DATA1_7  = p___constant_11x11xf32_5_5[7];
  assign \U312/DATA1_8  = p___constant_11x11xf32_5_5[8];
  assign \U312/DATA1_9  = p___constant_11x11xf32_5_5[9];
  assign \U312/DATA1_10  = p___constant_11x11xf32_5_5[10];
  assign \U312/DATA1_11  = p___constant_11x11xf32_5_5[11];
  assign \U307/DATA1_5  = p___constant_11x11xf32_5_6[5];
  assign \U307/DATA1_6  = p___constant_11x11xf32_5_6[6];
  assign \U307/DATA1_7  = p___constant_11x11xf32_5_6[7];
  assign \U307/DATA1_8  = p___constant_11x11xf32_5_6[8];
  assign \U307/DATA1_9  = p___constant_11x11xf32_5_6[9];
  assign \U307/DATA1_10  = p___constant_11x11xf32_5_6[10];
  assign \U307/DATA1_11  = p___constant_11x11xf32_5_6[11];
  assign \U302/DATA1_1  = p___constant_11x11xf32_5_7[1];
  assign \U302/DATA1_2  = p___constant_11x11xf32_5_7[2];
  assign \U302/DATA1_3  = p___constant_11x11xf32_5_7[3];
  assign \U302/DATA1_4  = p___constant_11x11xf32_5_7[4];
  assign \U302/DATA1_5  = p___constant_11x11xf32_5_7[5];
  assign \U302/DATA1_6  = p___constant_11x11xf32_5_7[6];
  assign \U302/DATA1_7  = p___constant_11x11xf32_5_7[7];
  assign \U302/DATA1_8  = p___constant_11x11xf32_5_7[8];
  assign \U302/DATA1_9  = p___constant_11x11xf32_5_7[9];
  assign \U302/DATA1_10  = p___constant_11x11xf32_5_7[10];
  assign \U302/DATA1_11  = p___constant_11x11xf32_5_7[11];
  assign \U297/DATA1_7  = p___constant_11x11xf32_5_8[7];
  assign \U297/DATA1_8  = p___constant_11x11xf32_5_8[8];
  assign \U297/DATA1_9  = p___constant_11x11xf32_5_8[9];
  assign \U297/DATA1_10  = p___constant_11x11xf32_5_8[10];
  assign \U297/DATA1_11  = p___constant_11x11xf32_5_8[11];
  assign \U292/DATA1_1  = p___constant_11x11xf32_5_9[1];
  assign \U292/DATA1_2  = p___constant_11x11xf32_5_9[2];
  assign \U292/DATA1_3  = p___constant_11x11xf32_5_9[3];
  assign \U292/DATA1_4  = p___constant_11x11xf32_5_9[4];
  assign \U292/DATA1_5  = p___constant_11x11xf32_5_9[5];
  assign \U292/DATA1_6  = p___constant_11x11xf32_5_9[6];
  assign \U292/DATA1_7  = p___constant_11x11xf32_5_9[7];
  assign \U292/DATA1_8  = p___constant_11x11xf32_5_9[8];
  assign \U292/DATA1_9  = p___constant_11x11xf32_5_9[9];
  assign \U292/DATA1_10  = p___constant_11x11xf32_5_9[10];
  assign \U292/DATA1_11  = p___constant_11x11xf32_5_9[11];
  assign \U287/DATA1_2  = p___constant_11x11xf32_5_10[2];
  assign \U287/DATA1_3  = p___constant_11x11xf32_5_10[3];
  assign \U287/DATA1_4  = p___constant_11x11xf32_5_10[4];
  assign \U287/DATA1_5  = p___constant_11x11xf32_5_10[5];
  assign \U287/DATA1_6  = p___constant_11x11xf32_5_10[6];
  assign \U287/DATA1_7  = p___constant_11x11xf32_5_10[7];
  assign \U287/DATA1_8  = p___constant_11x11xf32_5_10[8];
  assign \U287/DATA1_9  = p___constant_11x11xf32_5_10[9];
  assign \U287/DATA1_10  = p___constant_11x11xf32_5_10[10];
  assign \U287/DATA1_11  = p___constant_11x11xf32_5_10[11];
  assign \U282/DATA1_1  = p___constant_11xf32_5[1];
  assign \U282/DATA1_2  = p___constant_11xf32_5[2];
  assign \U282/DATA1_3  = p___constant_11xf32_5[3];
  assign \U282/DATA1_4  = p___constant_11xf32_5[4];
  assign \U282/DATA1_5  = p___constant_11xf32_5[5];
  assign \U282/DATA1_6  = p___constant_11xf32_5[6];
  assign \U282/DATA1_7  = p___constant_11xf32_5[7];
  assign \U282/DATA1_8  = p___constant_11xf32_5[8];
  assign \U282/DATA1_9  = p___constant_11xf32_5[9];
  assign \U282/DATA1_10  = p___constant_11xf32_5[10];
  assign \U282/DATA1_11  = p___constant_11xf32_5[11];
  assign \U279/DATA2_1  = p___constant_11x11xf32_6_0[1];
  assign \U279/DATA2_2  = p___constant_11x11xf32_6_0[2];
  assign \U279/DATA2_3  = p___constant_11x11xf32_6_0[3];
  assign \U279/DATA2_4  = p___constant_11x11xf32_6_0[4];
  assign \U279/DATA2_5  = p___constant_11x11xf32_6_0[5];
  assign \U279/DATA2_6  = p___constant_11x11xf32_6_0[6];
  assign \U279/DATA2_7  = p___constant_11x11xf32_6_0[7];
  assign \U279/DATA2_8  = p___constant_11x11xf32_6_0[8];
  assign \U279/DATA2_9  = p___constant_11x11xf32_6_0[9];
  assign \U279/DATA2_10  = p___constant_11x11xf32_6_0[10];
  assign \U279/DATA2_11  = p___constant_11x11xf32_6_0[11];
  assign \U279/DATA1_1  = p___constant_11x11xf32_6_1[1];
  assign \U279/DATA1_2  = p___constant_11x11xf32_6_1[2];
  assign \U279/DATA1_3  = p___constant_11x11xf32_6_1[3];
  assign \U279/DATA1_4  = p___constant_11x11xf32_6_1[4];
  assign \U279/DATA1_5  = p___constant_11x11xf32_6_1[5];
  assign \U279/DATA1_6  = p___constant_11x11xf32_6_1[6];
  assign \U279/DATA1_7  = p___constant_11x11xf32_6_1[7];
  assign \U279/DATA1_8  = p___constant_11x11xf32_6_1[8];
  assign \U279/DATA1_9  = p___constant_11x11xf32_6_1[9];
  assign \U279/DATA1_10  = p___constant_11x11xf32_6_1[10];
  assign \U279/DATA1_11  = p___constant_11x11xf32_6_1[11];
  assign \U274/DATA1_2  = p___constant_11x11xf32_6_2[2];
  assign \U274/DATA1_3  = p___constant_11x11xf32_6_2[3];
  assign \U274/DATA1_4  = p___constant_11x11xf32_6_2[4];
  assign \U274/DATA1_5  = p___constant_11x11xf32_6_2[5];
  assign \U274/DATA1_6  = p___constant_11x11xf32_6_2[6];
  assign \U274/DATA1_7  = p___constant_11x11xf32_6_2[7];
  assign \U274/DATA1_8  = p___constant_11x11xf32_6_2[8];
  assign \U274/DATA1_9  = p___constant_11x11xf32_6_2[9];
  assign \U274/DATA1_10  = p___constant_11x11xf32_6_2[10];
  assign \U274/DATA1_11  = p___constant_11x11xf32_6_2[11];
  assign \U269/DATA1_1  = p___constant_11x11xf32_6_3[1];
  assign \U269/DATA1_2  = p___constant_11x11xf32_6_3[2];
  assign \U269/DATA1_3  = p___constant_11x11xf32_6_3[3];
  assign \U269/DATA1_4  = p___constant_11x11xf32_6_3[4];
  assign \U269/DATA1_5  = p___constant_11x11xf32_6_3[5];
  assign \U269/DATA1_6  = p___constant_11x11xf32_6_3[6];
  assign \U269/DATA1_7  = p___constant_11x11xf32_6_3[7];
  assign \U269/DATA1_8  = p___constant_11x11xf32_6_3[8];
  assign \U269/DATA1_9  = p___constant_11x11xf32_6_3[9];
  assign \U269/DATA1_10  = p___constant_11x11xf32_6_3[10];
  assign \U269/DATA1_11  = p___constant_11x11xf32_6_3[11];
  assign \U264/DATA1_1  = p___constant_11x11xf32_6_4[1];
  assign \U264/DATA1_2  = p___constant_11x11xf32_6_4[2];
  assign \U264/DATA1_3  = p___constant_11x11xf32_6_4[3];
  assign \U264/DATA1_4  = p___constant_11x11xf32_6_4[4];
  assign \U264/DATA1_5  = p___constant_11x11xf32_6_4[5];
  assign \U264/DATA1_6  = p___constant_11x11xf32_6_4[6];
  assign \U264/DATA1_7  = p___constant_11x11xf32_6_4[7];
  assign \U264/DATA1_8  = p___constant_11x11xf32_6_4[8];
  assign \U264/DATA1_9  = p___constant_11x11xf32_6_4[9];
  assign \U264/DATA1_10  = p___constant_11x11xf32_6_4[10];
  assign \U264/DATA1_11  = p___constant_11x11xf32_6_4[11];
  assign \U254/DATA1_1  = p___constant_11x11xf32_6_6[1];
  assign \U254/DATA1_2  = p___constant_11x11xf32_6_6[2];
  assign \U254/DATA1_3  = p___constant_11x11xf32_6_6[3];
  assign \U254/DATA1_4  = p___constant_11x11xf32_6_6[4];
  assign \U254/DATA1_5  = p___constant_11x11xf32_6_6[5];
  assign \U254/DATA1_6  = p___constant_11x11xf32_6_6[6];
  assign \U254/DATA1_7  = p___constant_11x11xf32_6_6[7];
  assign \U254/DATA1_8  = p___constant_11x11xf32_6_6[8];
  assign \U254/DATA1_9  = p___constant_11x11xf32_6_6[9];
  assign \U254/DATA1_10  = p___constant_11x11xf32_6_6[10];
  assign \U254/DATA1_11  = p___constant_11x11xf32_6_6[11];
  assign \U249/DATA1_2  = p___constant_11x11xf32_6_7[2];
  assign \U249/DATA1_3  = p___constant_11x11xf32_6_7[3];
  assign \U249/DATA1_4  = p___constant_11x11xf32_6_7[4];
  assign \U249/DATA1_5  = p___constant_11x11xf32_6_7[5];
  assign \U249/DATA1_6  = p___constant_11x11xf32_6_7[6];
  assign \U249/DATA1_7  = p___constant_11x11xf32_6_7[7];
  assign \U249/DATA1_8  = p___constant_11x11xf32_6_7[8];
  assign \U249/DATA1_9  = p___constant_11x11xf32_6_7[9];
  assign \U249/DATA1_10  = p___constant_11x11xf32_6_7[10];
  assign \U249/DATA1_11  = p___constant_11x11xf32_6_7[11];
  assign \U244/DATA1_3  = p___constant_11x11xf32_6_8[3];
  assign \U244/DATA1_4  = p___constant_11x11xf32_6_8[4];
  assign \U244/DATA1_5  = p___constant_11x11xf32_6_8[5];
  assign \U244/DATA1_6  = p___constant_11x11xf32_6_8[6];
  assign \U244/DATA1_7  = p___constant_11x11xf32_6_8[7];
  assign \U244/DATA1_8  = p___constant_11x11xf32_6_8[8];
  assign \U244/DATA1_9  = p___constant_11x11xf32_6_8[9];
  assign \U244/DATA1_10  = p___constant_11x11xf32_6_8[10];
  assign \U244/DATA1_11  = p___constant_11x11xf32_6_8[11];
  assign \U239/DATA1_1  = p___constant_11x11xf32_6_9[1];
  assign \U239/DATA1_2  = p___constant_11x11xf32_6_9[2];
  assign \U239/DATA1_3  = p___constant_11x11xf32_6_9[3];
  assign \U239/DATA1_4  = p___constant_11x11xf32_6_9[4];
  assign \U239/DATA1_5  = p___constant_11x11xf32_6_9[5];
  assign \U239/DATA1_6  = p___constant_11x11xf32_6_9[6];
  assign \U239/DATA1_7  = p___constant_11x11xf32_6_9[7];
  assign \U239/DATA1_8  = p___constant_11x11xf32_6_9[8];
  assign \U239/DATA1_9  = p___constant_11x11xf32_6_9[9];
  assign \U239/DATA1_10  = p___constant_11x11xf32_6_9[10];
  assign \U239/DATA1_11  = p___constant_11x11xf32_6_9[11];
  assign \U234/DATA1_1  = p___constant_11x11xf32_6_10[1];
  assign \U234/DATA1_2  = p___constant_11x11xf32_6_10[2];
  assign \U234/DATA1_3  = p___constant_11x11xf32_6_10[3];
  assign \U234/DATA1_4  = p___constant_11x11xf32_6_10[4];
  assign \U234/DATA1_5  = p___constant_11x11xf32_6_10[5];
  assign \U234/DATA1_6  = p___constant_11x11xf32_6_10[6];
  assign \U234/DATA1_7  = p___constant_11x11xf32_6_10[7];
  assign \U234/DATA1_8  = p___constant_11x11xf32_6_10[8];
  assign \U234/DATA1_9  = p___constant_11x11xf32_6_10[9];
  assign \U234/DATA1_10  = p___constant_11x11xf32_6_10[10];
  assign \U234/DATA1_11  = p___constant_11x11xf32_6_10[11];
  assign \U229/DATA1_6  = p___constant_11xf32_6[6];
  assign \U229/DATA1_7  = p___constant_11xf32_6[7];
  assign \U229/DATA1_8  = p___constant_11xf32_6[8];
  assign \U229/DATA1_9  = p___constant_11xf32_6[9];
  assign \U229/DATA1_10  = p___constant_11xf32_6[10];
  assign \U229/DATA1_11  = p___constant_11xf32_6[11];
  assign \U223/DATA2_6  = p___constant_11x11xf32_7_0[6];
  assign \U223/DATA2_7  = p___constant_11x11xf32_7_0[7];
  assign \U223/DATA2_8  = p___constant_11x11xf32_7_0[8];
  assign \U223/DATA2_9  = p___constant_11x11xf32_7_0[9];
  assign \U223/DATA2_10  = p___constant_11x11xf32_7_0[10];
  assign \U223/DATA2_11  = p___constant_11x11xf32_7_0[11];
  assign \U223/DATA1_6  = p___constant_11x11xf32_7_1[6];
  assign \U223/DATA1_7  = p___constant_11x11xf32_7_1[7];
  assign \U223/DATA1_8  = p___constant_11x11xf32_7_1[8];
  assign \U223/DATA1_9  = p___constant_11x11xf32_7_1[9];
  assign \U223/DATA1_10  = p___constant_11x11xf32_7_1[10];
  assign \U223/DATA1_11  = p___constant_11x11xf32_7_1[11];
  assign \U218/DATA1_6  = p___constant_11x11xf32_7_2[6];
  assign \U218/DATA1_7  = p___constant_11x11xf32_7_2[7];
  assign \U218/DATA1_8  = p___constant_11x11xf32_7_2[8];
  assign \U218/DATA1_9  = p___constant_11x11xf32_7_2[9];
  assign \U218/DATA1_10  = p___constant_11x11xf32_7_2[10];
  assign \U218/DATA1_11  = p___constant_11x11xf32_7_2[11];
  assign \U213/DATA1_6  = p___constant_11x11xf32_7_3[6];
  assign \U213/DATA1_7  = p___constant_11x11xf32_7_3[7];
  assign \U213/DATA1_8  = p___constant_11x11xf32_7_3[8];
  assign \U213/DATA1_9  = p___constant_11x11xf32_7_3[9];
  assign \U213/DATA1_10  = p___constant_11x11xf32_7_3[10];
  assign \U213/DATA1_11  = p___constant_11x11xf32_7_3[11];
  assign \U208/DATA1_6  = p___constant_11x11xf32_7_4[6];
  assign \U208/DATA1_7  = p___constant_11x11xf32_7_4[7];
  assign \U208/DATA1_8  = p___constant_11x11xf32_7_4[8];
  assign \U208/DATA1_9  = p___constant_11x11xf32_7_4[9];
  assign \U208/DATA1_10  = p___constant_11x11xf32_7_4[10];
  assign \U208/DATA1_11  = p___constant_11x11xf32_7_4[11];
  assign \U203/DATA1_7  = p___constant_11x11xf32_7_5[7];
  assign \U203/DATA1_8  = p___constant_11x11xf32_7_5[8];
  assign \U203/DATA1_9  = p___constant_11x11xf32_7_5[9];
  assign \U203/DATA1_10  = p___constant_11x11xf32_7_5[10];
  assign \U203/DATA1_11  = p___constant_11x11xf32_7_5[11];
  assign \U198/DATA1_7  = p___constant_11x11xf32_7_6[7];
  assign \U198/DATA1_8  = p___constant_11x11xf32_7_6[8];
  assign \U198/DATA1_9  = p___constant_11x11xf32_7_6[9];
  assign \U198/DATA1_10  = p___constant_11x11xf32_7_6[10];
  assign \U198/DATA1_11  = p___constant_11x11xf32_7_6[11];
  assign \U193/DATA1_7  = p___constant_11x11xf32_7_7[7];
  assign \U193/DATA1_8  = p___constant_11x11xf32_7_7[8];
  assign \U193/DATA1_9  = p___constant_11x11xf32_7_7[9];
  assign \U193/DATA1_10  = p___constant_11x11xf32_7_7[10];
  assign \U193/DATA1_11  = p___constant_11x11xf32_7_7[11];
  assign \U188/DATA1_7  = p___constant_11x11xf32_7_8[7];
  assign \U188/DATA1_8  = p___constant_11x11xf32_7_8[8];
  assign \U188/DATA1_9  = p___constant_11x11xf32_7_8[9];
  assign \U188/DATA1_10  = p___constant_11x11xf32_7_8[10];
  assign \U188/DATA1_11  = p___constant_11x11xf32_7_8[11];
  assign \U183/DATA1_7  = p___constant_11x11xf32_7_9[7];
  assign \U183/DATA1_8  = p___constant_11x11xf32_7_9[8];
  assign \U183/DATA1_9  = p___constant_11x11xf32_7_9[9];
  assign \U183/DATA1_10  = p___constant_11x11xf32_7_9[10];
  assign \U183/DATA1_11  = p___constant_11x11xf32_7_9[11];
  assign \U178/DATA1_7  = p___constant_11x11xf32_7_10[7];
  assign \U178/DATA1_8  = p___constant_11x11xf32_7_10[8];
  assign \U178/DATA1_9  = p___constant_11x11xf32_7_10[9];
  assign \U178/DATA1_10  = p___constant_11x11xf32_7_10[10];
  assign \U178/DATA1_11  = p___constant_11x11xf32_7_10[11];
  assign \U173/DATA1_2  = p___constant_11xf32_7[2];
  assign \U173/DATA1_3  = p___constant_11xf32_7[3];
  assign \U173/DATA1_4  = p___constant_11xf32_7[4];
  assign \U173/DATA1_5  = p___constant_11xf32_7[5];
  assign \U173/DATA1_6  = p___constant_11xf32_7[6];
  assign \U173/DATA1_7  = p___constant_11xf32_7[7];
  assign \U173/DATA1_8  = p___constant_11xf32_7[8];
  assign \U173/DATA1_9  = p___constant_11xf32_7[9];
  assign \U173/DATA1_10  = p___constant_11xf32_7[10];
  assign \U173/DATA1_11  = p___constant_11xf32_7[11];
  assign \U170/DATA2_2  = p___constant_11x11xf32_8_0[2];
  assign \U170/DATA2_3  = p___constant_11x11xf32_8_0[3];
  assign \U170/DATA2_4  = p___constant_11x11xf32_8_0[4];
  assign \U170/DATA2_5  = p___constant_11x11xf32_8_0[5];
  assign \U170/DATA2_6  = p___constant_11x11xf32_8_0[6];
  assign \U170/DATA2_7  = p___constant_11x11xf32_8_0[7];
  assign \U170/DATA2_8  = p___constant_11x11xf32_8_0[8];
  assign \U170/DATA2_9  = p___constant_11x11xf32_8_0[9];
  assign \U170/DATA2_10  = p___constant_11x11xf32_8_0[10];
  assign \U170/DATA2_11  = p___constant_11x11xf32_8_0[11];
  assign \U170/DATA1_2  = p___constant_11x11xf32_8_1[2];
  assign \U170/DATA1_3  = p___constant_11x11xf32_8_1[3];
  assign \U170/DATA1_4  = p___constant_11x11xf32_8_1[4];
  assign \U170/DATA1_5  = p___constant_11x11xf32_8_1[5];
  assign \U170/DATA1_6  = p___constant_11x11xf32_8_1[6];
  assign \U170/DATA1_7  = p___constant_11x11xf32_8_1[7];
  assign \U170/DATA1_8  = p___constant_11x11xf32_8_1[8];
  assign \U170/DATA1_9  = p___constant_11x11xf32_8_1[9];
  assign \U170/DATA1_10  = p___constant_11x11xf32_8_1[10];
  assign \U170/DATA1_11  = p___constant_11x11xf32_8_1[11];
  assign \U165/DATA1_2  = p___constant_11x11xf32_8_2[2];
  assign \U165/DATA1_3  = p___constant_11x11xf32_8_2[3];
  assign \U165/DATA1_4  = p___constant_11x11xf32_8_2[4];
  assign \U165/DATA1_5  = p___constant_11x11xf32_8_2[5];
  assign \U165/DATA1_6  = p___constant_11x11xf32_8_2[6];
  assign \U165/DATA1_7  = p___constant_11x11xf32_8_2[7];
  assign \U165/DATA1_8  = p___constant_11x11xf32_8_2[8];
  assign \U165/DATA1_9  = p___constant_11x11xf32_8_2[9];
  assign \U165/DATA1_10  = p___constant_11x11xf32_8_2[10];
  assign \U165/DATA1_11  = p___constant_11x11xf32_8_2[11];
  assign \U160/DATA1_2  = p___constant_11x11xf32_8_3[2];
  assign \U160/DATA1_3  = p___constant_11x11xf32_8_3[3];
  assign \U160/DATA1_4  = p___constant_11x11xf32_8_3[4];
  assign \U160/DATA1_5  = p___constant_11x11xf32_8_3[5];
  assign \U160/DATA1_6  = p___constant_11x11xf32_8_3[6];
  assign \U160/DATA1_7  = p___constant_11x11xf32_8_3[7];
  assign \U160/DATA1_8  = p___constant_11x11xf32_8_3[8];
  assign \U160/DATA1_9  = p___constant_11x11xf32_8_3[9];
  assign \U160/DATA1_10  = p___constant_11x11xf32_8_3[10];
  assign \U160/DATA1_11  = p___constant_11x11xf32_8_3[11];
  assign \U155/DATA1_2  = p___constant_11x11xf32_8_4[2];
  assign \U155/DATA1_3  = p___constant_11x11xf32_8_4[3];
  assign \U155/DATA1_4  = p___constant_11x11xf32_8_4[4];
  assign \U155/DATA1_5  = p___constant_11x11xf32_8_4[5];
  assign \U155/DATA1_6  = p___constant_11x11xf32_8_4[6];
  assign \U155/DATA1_7  = p___constant_11x11xf32_8_4[7];
  assign \U155/DATA1_8  = p___constant_11x11xf32_8_4[8];
  assign \U155/DATA1_9  = p___constant_11x11xf32_8_4[9];
  assign \U155/DATA1_10  = p___constant_11x11xf32_8_4[10];
  assign \U155/DATA1_11  = p___constant_11x11xf32_8_4[11];
  assign \U150/DATA1_2  = p___constant_11x11xf32_8_5[2];
  assign \U150/DATA1_3  = p___constant_11x11xf32_8_5[3];
  assign \U150/DATA1_4  = p___constant_11x11xf32_8_5[4];
  assign \U150/DATA1_5  = p___constant_11x11xf32_8_5[5];
  assign \U150/DATA1_6  = p___constant_11x11xf32_8_5[6];
  assign \U150/DATA1_7  = p___constant_11x11xf32_8_5[7];
  assign \U150/DATA1_8  = p___constant_11x11xf32_8_5[8];
  assign \U150/DATA1_9  = p___constant_11x11xf32_8_5[9];
  assign \U150/DATA1_10  = p___constant_11x11xf32_8_5[10];
  assign \U150/DATA1_11  = p___constant_11x11xf32_8_5[11];
  assign \U145/DATA1_2  = p___constant_11x11xf32_8_6[2];
  assign \U145/DATA1_3  = p___constant_11x11xf32_8_6[3];
  assign \U145/DATA1_4  = p___constant_11x11xf32_8_6[4];
  assign \U145/DATA1_5  = p___constant_11x11xf32_8_6[5];
  assign \U145/DATA1_6  = p___constant_11x11xf32_8_6[6];
  assign \U145/DATA1_7  = p___constant_11x11xf32_8_6[7];
  assign \U145/DATA1_8  = p___constant_11x11xf32_8_6[8];
  assign \U145/DATA1_9  = p___constant_11x11xf32_8_6[9];
  assign \U145/DATA1_10  = p___constant_11x11xf32_8_6[10];
  assign \U145/DATA1_11  = p___constant_11x11xf32_8_6[11];
  assign \U140/DATA1_0  = p___constant_11x11xf32_8_7[0];
  assign \U140/DATA1_1  = p___constant_11x11xf32_8_7[1];
  assign \U140/DATA1_2  = p___constant_11x11xf32_8_7[2];
  assign \U140/DATA1_3  = p___constant_11x11xf32_8_7[3];
  assign \U140/DATA1_4  = p___constant_11x11xf32_8_7[4];
  assign \U140/DATA1_5  = p___constant_11x11xf32_8_7[5];
  assign \U140/DATA1_6  = p___constant_11x11xf32_8_7[6];
  assign \U140/DATA1_7  = p___constant_11x11xf32_8_7[7];
  assign \U140/DATA1_8  = p___constant_11x11xf32_8_7[8];
  assign \U140/DATA1_9  = p___constant_11x11xf32_8_7[9];
  assign \U140/DATA1_10  = p___constant_11x11xf32_8_7[10];
  assign \U140/DATA1_11  = p___constant_11x11xf32_8_7[11];
  assign \U135/DATA1_0  = p___constant_11x11xf32_8_8[0];
  assign \U135/DATA1_1  = p___constant_11x11xf32_8_8[1];
  assign \U135/DATA1_2  = p___constant_11x11xf32_8_8[2];
  assign \U135/DATA1_3  = p___constant_11x11xf32_8_8[3];
  assign \U135/DATA1_4  = p___constant_11x11xf32_8_8[4];
  assign \U135/DATA1_5  = p___constant_11x11xf32_8_8[5];
  assign \U135/DATA1_6  = p___constant_11x11xf32_8_8[6];
  assign \U135/DATA1_7  = p___constant_11x11xf32_8_8[7];
  assign \U135/DATA1_8  = p___constant_11x11xf32_8_8[8];
  assign \U135/DATA1_9  = p___constant_11x11xf32_8_8[9];
  assign \U135/DATA1_10  = p___constant_11x11xf32_8_8[10];
  assign \U135/DATA1_11  = p___constant_11x11xf32_8_8[11];
  assign \U130/DATA1_0  = p___constant_11x11xf32_8_9[0];
  assign \U130/DATA1_1  = p___constant_11x11xf32_8_9[1];
  assign \U130/DATA1_2  = p___constant_11x11xf32_8_9[2];
  assign \U130/DATA1_3  = p___constant_11x11xf32_8_9[3];
  assign \U130/DATA1_4  = p___constant_11x11xf32_8_9[4];
  assign \U130/DATA1_5  = p___constant_11x11xf32_8_9[5];
  assign \U130/DATA1_6  = p___constant_11x11xf32_8_9[6];
  assign \U130/DATA1_7  = p___constant_11x11xf32_8_9[7];
  assign \U130/DATA1_8  = p___constant_11x11xf32_8_9[8];
  assign \U130/DATA1_9  = p___constant_11x11xf32_8_9[9];
  assign \U130/DATA1_10  = p___constant_11x11xf32_8_9[10];
  assign \U130/DATA1_11  = p___constant_11x11xf32_8_9[11];
  assign \U125/DATA1_0  = p___constant_11x11xf32_8_10[0];
  assign \U125/DATA1_1  = p___constant_11x11xf32_8_10[1];
  assign \U125/DATA1_2  = p___constant_11x11xf32_8_10[2];
  assign \U125/DATA1_3  = p___constant_11x11xf32_8_10[3];
  assign \U125/DATA1_4  = p___constant_11x11xf32_8_10[4];
  assign \U125/DATA1_5  = p___constant_11x11xf32_8_10[5];
  assign \U125/DATA1_6  = p___constant_11x11xf32_8_10[6];
  assign \U125/DATA1_7  = p___constant_11x11xf32_8_10[7];
  assign \U125/DATA1_8  = p___constant_11x11xf32_8_10[8];
  assign \U125/DATA1_9  = p___constant_11x11xf32_8_10[9];
  assign \U125/DATA1_10  = p___constant_11x11xf32_8_10[10];
  assign \U125/DATA1_11  = p___constant_11x11xf32_8_10[11];
  assign \U120/DATA1_0  = p___constant_11xf32_8[0];
  assign \U120/DATA1_1  = p___constant_11xf32_8[1];
  assign \U120/DATA1_2  = p___constant_11xf32_8[2];
  assign \U120/DATA1_3  = p___constant_11xf32_8[3];
  assign \U120/DATA1_4  = p___constant_11xf32_8[4];
  assign \U120/DATA1_5  = p___constant_11xf32_8[5];
  assign \U120/DATA1_6  = p___constant_11xf32_8[6];
  assign \U120/DATA1_7  = p___constant_11xf32_8[7];
  assign \U120/DATA1_8  = p___constant_11xf32_8[8];
  assign \U120/DATA1_9  = p___constant_11xf32_8[9];
  assign \U120/DATA1_10  = p___constant_11xf32_8[10];
  assign \U120/DATA1_11  = p___constant_11xf32_8[11];
  assign \U108/DATA2_0  = p___constant_11x11xf32_9_0[0];
  assign \U108/DATA2_1  = p___constant_11x11xf32_9_0[1];
  assign \U108/DATA2_2  = p___constant_11x11xf32_9_0[2];
  assign \U108/DATA2_3  = p___constant_11x11xf32_9_0[3];
  assign \U108/DATA2_4  = p___constant_11x11xf32_9_0[4];
  assign \U108/DATA2_5  = p___constant_11x11xf32_9_0[5];
  assign \U108/DATA2_6  = p___constant_11x11xf32_9_0[6];
  assign \U108/DATA2_7  = p___constant_11x11xf32_9_0[7];
  assign \U108/DATA2_8  = p___constant_11x11xf32_9_0[8];
  assign \U108/DATA2_9  = p___constant_11x11xf32_9_0[9];
  assign \U108/DATA2_10  = p___constant_11x11xf32_9_0[10];
  assign \U108/DATA2_11  = p___constant_11x11xf32_9_0[11];
  assign \U108/DATA1_0  = p___constant_11x11xf32_9_1[0];
  assign \U108/DATA1_1  = p___constant_11x11xf32_9_1[1];
  assign \U108/DATA1_2  = p___constant_11x11xf32_9_1[2];
  assign \U108/DATA1_3  = p___constant_11x11xf32_9_1[3];
  assign \U108/DATA1_4  = p___constant_11x11xf32_9_1[4];
  assign \U108/DATA1_5  = p___constant_11x11xf32_9_1[5];
  assign \U108/DATA1_6  = p___constant_11x11xf32_9_1[6];
  assign \U108/DATA1_7  = p___constant_11x11xf32_9_1[7];
  assign \U108/DATA1_8  = p___constant_11x11xf32_9_1[8];
  assign \U108/DATA1_9  = p___constant_11x11xf32_9_1[9];
  assign \U108/DATA1_10  = p___constant_11x11xf32_9_1[10];
  assign \U108/DATA1_11  = p___constant_11x11xf32_9_1[11];
  assign \U103/DATA1_0  = p___constant_11x11xf32_9_2[0];
  assign \U103/DATA1_1  = p___constant_11x11xf32_9_2[1];
  assign \U103/DATA1_2  = p___constant_11x11xf32_9_2[2];
  assign \U103/DATA1_3  = p___constant_11x11xf32_9_2[3];
  assign \U103/DATA1_4  = p___constant_11x11xf32_9_2[4];
  assign \U103/DATA1_5  = p___constant_11x11xf32_9_2[5];
  assign \U103/DATA1_6  = p___constant_11x11xf32_9_2[6];
  assign \U103/DATA1_7  = p___constant_11x11xf32_9_2[7];
  assign \U103/DATA1_8  = p___constant_11x11xf32_9_2[8];
  assign \U103/DATA1_9  = p___constant_11x11xf32_9_2[9];
  assign \U103/DATA1_10  = p___constant_11x11xf32_9_2[10];
  assign \U103/DATA1_11  = p___constant_11x11xf32_9_2[11];
  assign \U98/DATA1_0  = p___constant_11x11xf32_9_3[0];
  assign \U98/DATA1_1  = p___constant_11x11xf32_9_3[1];
  assign \U98/DATA1_2  = p___constant_11x11xf32_9_3[2];
  assign \U98/DATA1_3  = p___constant_11x11xf32_9_3[3];
  assign \U98/DATA1_4  = p___constant_11x11xf32_9_3[4];
  assign \U98/DATA1_5  = p___constant_11x11xf32_9_3[5];
  assign \U98/DATA1_6  = p___constant_11x11xf32_9_3[6];
  assign \U98/DATA1_7  = p___constant_11x11xf32_9_3[7];
  assign \U98/DATA1_8  = p___constant_11x11xf32_9_3[8];
  assign \U98/DATA1_9  = p___constant_11x11xf32_9_3[9];
  assign \U98/DATA1_10  = p___constant_11x11xf32_9_3[10];
  assign \U98/DATA1_11  = p___constant_11x11xf32_9_3[11];
  assign \U93/DATA1_5  = p___constant_11x11xf32_9_4[5];
  assign \U93/DATA1_6  = p___constant_11x11xf32_9_4[6];
  assign \U93/DATA1_7  = p___constant_11x11xf32_9_4[7];
  assign \U93/DATA1_8  = p___constant_11x11xf32_9_4[8];
  assign \U93/DATA1_9  = p___constant_11x11xf32_9_4[9];
  assign \U93/DATA1_10  = p___constant_11x11xf32_9_4[10];
  assign \U93/DATA1_11  = p___constant_11x11xf32_9_4[11];
  assign \U88/DATA1_1  = p___constant_11x11xf32_9_5[1];
  assign \U88/DATA1_2  = p___constant_11x11xf32_9_5[2];
  assign \U88/DATA1_3  = p___constant_11x11xf32_9_5[3];
  assign \U88/DATA1_4  = p___constant_11x11xf32_9_5[4];
  assign \U88/DATA1_5  = p___constant_11x11xf32_9_5[5];
  assign \U88/DATA1_6  = p___constant_11x11xf32_9_5[6];
  assign \U88/DATA1_7  = p___constant_11x11xf32_9_5[7];
  assign \U88/DATA1_8  = p___constant_11x11xf32_9_5[8];
  assign \U88/DATA1_9  = p___constant_11x11xf32_9_5[9];
  assign \U88/DATA1_10  = p___constant_11x11xf32_9_5[10];
  assign \U88/DATA1_11  = p___constant_11x11xf32_9_5[11];
  assign \U83/DATA1_4  = p___constant_11x11xf32_9_6[4];
  assign \U83/DATA1_5  = p___constant_11x11xf32_9_6[5];
  assign \U83/DATA1_6  = p___constant_11x11xf32_9_6[6];
  assign \U83/DATA1_7  = p___constant_11x11xf32_9_6[7];
  assign \U83/DATA1_8  = p___constant_11x11xf32_9_6[8];
  assign \U83/DATA1_9  = p___constant_11x11xf32_9_6[9];
  assign \U83/DATA1_10  = p___constant_11x11xf32_9_6[10];
  assign \U83/DATA1_11  = p___constant_11x11xf32_9_6[11];
  assign \U78/DATA1_9  = p___constant_11x11xf32_9_7[9];
  assign \U78/DATA1_10  = p___constant_11x11xf32_9_7[10];
  assign \U78/DATA1_11  = p___constant_11x11xf32_9_7[11];
  assign \U73/DATA1_1  = p___constant_11x11xf32_9_8[1];
  assign \U73/DATA1_2  = p___constant_11x11xf32_9_8[2];
  assign \U73/DATA1_3  = p___constant_11x11xf32_9_8[3];
  assign \U73/DATA1_4  = p___constant_11x11xf32_9_8[4];
  assign \U73/DATA1_5  = p___constant_11x11xf32_9_8[5];
  assign \U73/DATA1_6  = p___constant_11x11xf32_9_8[6];
  assign \U73/DATA1_7  = p___constant_11x11xf32_9_8[7];
  assign \U73/DATA1_8  = p___constant_11x11xf32_9_8[8];
  assign \U73/DATA1_9  = p___constant_11x11xf32_9_8[9];
  assign \U73/DATA1_10  = p___constant_11x11xf32_9_8[10];
  assign \U73/DATA1_11  = p___constant_11x11xf32_9_8[11];
  assign \U68/DATA1_6  = p___constant_11x11xf32_9_9[6];
  assign \U68/DATA1_7  = p___constant_11x11xf32_9_9[7];
  assign \U68/DATA1_8  = p___constant_11x11xf32_9_9[8];
  assign \U68/DATA1_9  = p___constant_11x11xf32_9_9[9];
  assign \U68/DATA1_10  = p___constant_11x11xf32_9_9[10];
  assign \U68/DATA1_11  = p___constant_11x11xf32_9_9[11];
  assign \U63/DATA1_11  = p___constant_11x11xf32_9_10[11];
  assign \U58/DATA1_4  = p___constant_11xf32_9[4];
  assign \U58/DATA1_5  = p___constant_11xf32_9[5];
  assign \U58/DATA1_6  = p___constant_11xf32_9[6];
  assign \U58/DATA1_7  = p___constant_11xf32_9[7];
  assign \U58/DATA1_8  = p___constant_11xf32_9[8];
  assign \U58/DATA1_9  = p___constant_11xf32_9[9];
  assign \U58/DATA1_10  = p___constant_11xf32_9[10];
  assign \U58/DATA1_11  = p___constant_11xf32_9[11];
  assign \U55/DATA2_11  = p___constant_11x11xf32_10_0[11];
  assign \U55/DATA1_11  = p___constant_11x11xf32_10_1[11];
  assign \U50/DATA1_4  = p___constant_11x11xf32_10_2[4];
  assign \U50/DATA1_5  = p___constant_11x11xf32_10_2[5];
  assign \U50/DATA1_6  = p___constant_11x11xf32_10_2[6];
  assign \U50/DATA1_7  = p___constant_11x11xf32_10_2[7];
  assign \U50/DATA1_8  = p___constant_11x11xf32_10_2[8];
  assign \U50/DATA1_9  = p___constant_11x11xf32_10_2[9];
  assign \U50/DATA1_10  = p___constant_11x11xf32_10_2[10];
  assign \U50/DATA1_11  = p___constant_11x11xf32_10_2[11];
  assign \U45/DATA1_5  = p___constant_11x11xf32_10_3[5];
  assign \U45/DATA1_6  = p___constant_11x11xf32_10_3[6];
  assign \U45/DATA1_7  = p___constant_11x11xf32_10_3[7];
  assign \U45/DATA1_8  = p___constant_11x11xf32_10_3[8];
  assign \U45/DATA1_9  = p___constant_11x11xf32_10_3[9];
  assign \U45/DATA1_10  = p___constant_11x11xf32_10_3[10];
  assign \U45/DATA1_11  = p___constant_11x11xf32_10_3[11];
  assign \U40/DATA1_1  = p___constant_11x11xf32_10_4[1];
  assign \U40/DATA1_2  = p___constant_11x11xf32_10_4[2];
  assign \U40/DATA1_3  = p___constant_11x11xf32_10_4[3];
  assign \U40/DATA1_4  = p___constant_11x11xf32_10_4[4];
  assign \U40/DATA1_5  = p___constant_11x11xf32_10_4[5];
  assign \U40/DATA1_6  = p___constant_11x11xf32_10_4[6];
  assign \U40/DATA1_7  = p___constant_11x11xf32_10_4[7];
  assign \U40/DATA1_8  = p___constant_11x11xf32_10_4[8];
  assign \U40/DATA1_9  = p___constant_11x11xf32_10_4[9];
  assign \U40/DATA1_10  = p___constant_11x11xf32_10_4[10];
  assign \U40/DATA1_11  = p___constant_11x11xf32_10_4[11];
  assign \U35/DATA1_4  = p___constant_11x11xf32_10_5[4];
  assign \U35/DATA1_5  = p___constant_11x11xf32_10_5[5];
  assign \U35/DATA1_6  = p___constant_11x11xf32_10_5[6];
  assign \U35/DATA1_7  = p___constant_11x11xf32_10_5[7];
  assign \U35/DATA1_8  = p___constant_11x11xf32_10_5[8];
  assign \U35/DATA1_9  = p___constant_11x11xf32_10_5[9];
  assign \U35/DATA1_10  = p___constant_11x11xf32_10_5[10];
  assign \U35/DATA1_11  = p___constant_11x11xf32_10_5[11];
  assign \U30/DATA1_9  = p___constant_11x11xf32_10_6[9];
  assign \U30/DATA1_10  = p___constant_11x11xf32_10_6[10];
  assign \U30/DATA1_11  = p___constant_11x11xf32_10_6[11];
  assign \U25/DATA1_1  = p___constant_11x11xf32_10_7[1];
  assign \U25/DATA1_2  = p___constant_11x11xf32_10_7[2];
  assign \U25/DATA1_3  = p___constant_11x11xf32_10_7[3];
  assign \U25/DATA1_4  = p___constant_11x11xf32_10_7[4];
  assign \U25/DATA1_5  = p___constant_11x11xf32_10_7[5];
  assign \U25/DATA1_6  = p___constant_11x11xf32_10_7[6];
  assign \U25/DATA1_7  = p___constant_11x11xf32_10_7[7];
  assign \U25/DATA1_8  = p___constant_11x11xf32_10_7[8];
  assign \U25/DATA1_9  = p___constant_11x11xf32_10_7[9];
  assign \U25/DATA1_10  = p___constant_11x11xf32_10_7[10];
  assign \U25/DATA1_11  = p___constant_11x11xf32_10_7[11];
  assign \U20/DATA1_6  = p___constant_11x11xf32_10_8[6];
  assign \U20/DATA1_7  = p___constant_11x11xf32_10_8[7];
  assign \U20/DATA1_8  = p___constant_11x11xf32_10_8[8];
  assign \U20/DATA1_9  = p___constant_11x11xf32_10_8[9];
  assign \U20/DATA1_10  = p___constant_11x11xf32_10_8[10];
  assign \U20/DATA1_11  = p___constant_11x11xf32_10_8[11];
  assign \U15/DATA1_11  = p___constant_11x11xf32_10_9[11];
  assign \U10/DATA1_9  = p___constant_11x11xf32_10_10[9];
  assign \U10/DATA1_10  = p___constant_11x11xf32_10_10[10];
  assign \U10/DATA1_11  = p___constant_11x11xf32_10_10[11];
  assign \U5/DATA1_9  = p___constant_11xf32_10[9];
  assign \U5/DATA1_10  = p___constant_11xf32_10[10];
  assign \U5/DATA1_11  = p___constant_11xf32_10[11];

  FADDX1 \fmul_0_0_0_0_10/add_2_root_add_321/U1_4  ( .A(
        \fmul_0_0_0_0_10/add_2_root_add_321/A[4] ), .B(
        \fmul_0_0_0_0_10/add_2_root_add_321/B[4] ), .CI(
        \fmul_0_0_0_0_10/add_2_root_add_321/carry[4] ), .CO(
        \fmul_0_0_0_0_10/add_2_root_add_321/carry[5] ), .S(
        \fmul_0_0_0_0_10/sub_1_root_add_321/A[4] ) );
  FADDX1 \fmul_0_0_0_0_10/add_2_root_add_321/U1_3  ( .A(
        \fmul_0_0_0_0_10/add_2_root_add_321/A[3] ), .B(
        \fmul_0_0_0_0_10/add_2_root_add_321/B[3] ), .CI(
        \fmul_0_0_0_0_10/add_2_root_add_321/carry[3] ), .CO(
        \fmul_0_0_0_0_10/add_2_root_add_321/carry[4] ), .S(
        \fmul_0_0_0_0_10/sub_1_root_add_321/A[3] ) );
  FADDX1 \fmul_0_0_0_0_10/add_2_root_add_321/U1_2  ( .A(
        \fmul_0_0_0_0_10/add_2_root_add_321/A[2] ), .B(
        \fmul_0_0_0_0_10/add_2_root_add_321/B[2] ), .CI(
        \fmul_0_0_0_0_10/add_2_root_add_321/carry[2] ), .CO(
        \fmul_0_0_0_0_10/add_2_root_add_321/carry[3] ), .S(
        \fmul_0_0_0_0_10/sub_1_root_add_321/A[2] ) );
  FADDX1 \fmul_0_0_0_0_10/add_2_root_add_321/U1_1  ( .A(
        \fmul_0_0_0_0_10/add_2_root_add_321/A[1] ), .B(
        \fmul_0_0_0_0_10/add_2_root_add_321/B[1] ), .CI(
        \fmul_0_0_0_0_10/add_2_root_add_321/carry[1] ), .CO(
        \fmul_0_0_0_0_10/add_2_root_add_321/carry[2] ), .S(
        \fmul_0_0_0_0_10/sub_1_root_add_321/A[1] ) );
  FADDX1 \fmul_0_0_0_0_10/add_2_root_add_321/U1_0  ( .A(
        \fmul_0_0_0_0_10/add_2_root_add_321/A[0] ), .B(
        \fmul_0_0_0_0_10/add_2_root_add_321/B[0] ), .CI(n14920), .CO(
        \fmul_0_0_0_0_10/add_2_root_add_321/carry[1] ), .S(
        \fmul_0_0_0_0_10/sub_1_root_add_321/A[0] ) );
  FADDX1 \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/U1_5  ( 
        .A(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/A[5] ), .B(\fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/B[5] ), 
        .CI(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/carry[5] ), .CO(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/carry[6] ), .S(\fadd_0_0_0_0_10/U21/DATA2_2 ) );
  FADDX1 \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/U1_4  ( 
        .A(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/A[4] ), .B(\fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/B[4] ), 
        .CI(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/carry[4] ), .CO(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/carry[5] ), .S(\fadd_0_0_0_0_10/U22/DATA1_3 ) );
  FADDX1 \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/U1_3  ( 
        .A(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/A[3] ), .B(\fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/B[3] ), 
        .CI(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/carry[3] ), .CO(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/carry[4] ), .S(\fadd_0_0_0_0_10/U22/DATA1_2 ) );
  FADDX1 \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/U1_2  ( 
        .A(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/A[2] ), .B(\fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/B[2] ), 
        .CI(n14138), .CO(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/carry[3] ), .S(\fadd_0_0_0_0_10/U22/DATA1_1 ) );
  FADDX1 \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_dualsubclose/sub_1_root_add_303/U2_4  ( 
        .A(n12794), .B(n14972), .CI(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_dualsubclose/sub_1_root_add_303/carry[4] ), .CO(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_dualsubclose/sub_1_root_add_303/carry[5] ), .S(\fadd_0_0_0_0_10/U24/DATA2_4 ) );
  FADDX1 \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_dualsubclose/sub_1_root_add_303/U2_3  ( 
        .A(\fadd_0_0_0_0_10/U25/Z_3 ), .B(n14969), .CI(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_dualsubclose/sub_1_root_add_303/carry[3] ), .CO(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_dualsubclose/sub_1_root_add_303/carry[4] ), .S(\fadd_0_0_0_0_10/U24/DATA2_3 ) );
  FADDX1 \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_dualsubclose/sub_1_root_add_303/U2_2  ( 
        .A(\fadd_0_0_0_0_10/U25/Z_2 ), .B(n14966), .CI(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_dualsubclose/sub_1_root_add_303/carry[2] ), .CO(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_dualsubclose/sub_1_root_add_303/carry[3] ), .S(\fadd_0_0_0_0_10/U24/DATA2_2 ) );
  FADDX1 \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_dualsubclose/sub_1_root_add_300/U2_3  ( 
        .A(\fadd_0_0_0_0_10/U29/Z_2 ), .B(n14970), .CI(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_dualsubclose/sub_1_root_add_300/carry[3] ), .CO(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_dualsubclose/sub_1_root_add_300/carry[4] ), .S(\fadd_0_0_0_0_10/U24/DATA1_3 ) );
  FADDX1 \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_dualsubclose/sub_1_root_add_300/U2_2  ( 
        .A(\fadd_0_0_0_0_10/U29/Z_1 ), .B(n14967), .CI(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_dualsubclose/sub_1_root_add_300/carry[2] ), .CO(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_dualsubclose/sub_1_root_add_300/carry[3] ), .S(\fadd_0_0_0_0_10/U24/DATA1_2 ) );
  FADDX1 \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_dualsubclose/sub_1_root_add_300/U2_1  ( 
        .A(\fadd_0_0_0_0_10/U29/Z_0 ), .B(n13467), .CI(n13401), .CO(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_dualsubclose/sub_1_root_add_300/carry[2] ), .S(\fadd_0_0_0_0_10/U24/DATA1_1 ) );
  FADDX1 \fadd_0_0_0_0_10/sub_784/U2_2  ( .A(\fadd_0_0_0_0_10/sub_784/A[2] ), 
        .B(n12871), .CI(\fadd_0_0_0_0_10/sub_784/carry[2] ), .CO(
        \fadd_0_0_0_0_10/sub_784/carry[3] ), .S(
        \fadd_0_0_0_0_10/sub_784/DIFF[2] ) );
  FADDX1 \fadd_0_0_0_0_10/sub_784/U2_1  ( .A(\fadd_0_0_0_0_10/sub_784/A[1] ), 
        .B(n12870), .CI(\fadd_0_0_0_0_10/sub_784/carry[1] ), .CO(
        \fadd_0_0_0_0_10/sub_784/carry[2] ), .S(
        \fadd_0_0_0_0_10/sub_784/DIFF[1] ) );
  FADDX1 \fadd_0_0_0_0_10/sub_710/U2_4  ( .A(n14983), .B(n12803), .CI(
        \fadd_0_0_0_0_10/sub_710/carry[4] ), .S(\fadd_0_0_0_0_10/U5/DATA1_4 )
         );
  FADDX1 \fadd_0_0_0_0_10/sub_710/U2_3  ( .A(n14982), .B(n12804), .CI(
        \fadd_0_0_0_0_10/sub_710/carry[3] ), .CO(
        \fadd_0_0_0_0_10/sub_710/carry[4] ), .S(\fadd_0_0_0_0_10/U5/DATA1_3 )
         );
  FADDX1 \fadd_0_0_0_0_10/sub_710/U2_2  ( .A(n14981), .B(n12805), .CI(
        \fadd_0_0_0_0_10/sub_710/carry[2] ), .CO(
        \fadd_0_0_0_0_10/sub_710/carry[3] ), .S(\fadd_0_0_0_0_10/U5/DATA1_2 )
         );
  FADDX1 \fadd_0_0_0_0_10/sub_710/U2_1  ( .A(n14980), .B(n12806), .CI(
        \fadd_0_0_0_0_10/sub_710/carry[1] ), .CO(
        \fadd_0_0_0_0_10/sub_710/carry[2] ), .S(\fadd_0_0_0_0_10/U5/DATA1_1 )
         );
  FADDX1 \fadd_0_0_0_0_10/sub_707/U2_4  ( .A(n14999), .B(n12810), .CI(
        \fadd_0_0_0_0_10/sub_707/carry[4] ), .CO(
        \fadd_0_0_0_0_10/sub_707/carry[5] ), .S(\fadd_0_0_0_0_10/U5/DATA2_4 )
         );
  FADDX1 \fadd_0_0_0_0_10/sub_707/U2_3  ( .A(n14998), .B(n12811), .CI(
        \fadd_0_0_0_0_10/sub_707/carry[3] ), .CO(
        \fadd_0_0_0_0_10/sub_707/carry[4] ), .S(\fadd_0_0_0_0_10/U5/DATA2_3 )
         );
  FADDX1 \fadd_0_0_0_0_10/sub_707/U2_2  ( .A(n14997), .B(n12812), .CI(
        \fadd_0_0_0_0_10/sub_707/carry[2] ), .CO(
        \fadd_0_0_0_0_10/sub_707/carry[3] ), .S(\fadd_0_0_0_0_10/U5/DATA2_2 )
         );
  FADDX1 \fadd_0_0_0_0_10/sub_707/U2_1  ( .A(n14996), .B(n12813), .CI(
        \fadd_0_0_0_0_10/sub_707/carry[1] ), .CO(
        \fadd_0_0_0_0_10/sub_707/carry[2] ), .S(\fadd_0_0_0_0_10/U5/DATA2_1 )
         );
  DFFX1 \current_fsm_reg[0]  ( .D(n13443), .CLK(clk), .QN(n13715) );
  DFFX1 \current_fsm_reg[1]  ( .D(n13442), .CLK(clk), .QN(n11608) );
  DFFX1 \current_fsm_reg[2]  ( .D(n13441), .CLK(clk), .QN(n11937) );
  DFFX1 \current_fsm_reg[3]  ( .D(n13440), .CLK(clk), .Q(n13674), .QN(n12837)
         );
  DFFX1 \current_fsm_reg[4]  ( .D(n13439), .CLK(clk), .QN(n11610) );
  DFFX1 \current_fsm_reg[5]  ( .D(n13438), .CLK(clk), .QN(n13631) );
  DFFX1 \current_fsm_reg[6]  ( .D(n13437), .CLK(clk), .Q(n13537), .QN(n12836)
         );
  DFFX1 \current_fsm_reg[7]  ( .D(n13436), .CLK(clk), .QN(n11611) );
  DFFX1 \current_fsm_reg[8]  ( .D(n13435), .CLK(clk), .QN(n13476) );
  DFFX1 \current_fsm_reg[9]  ( .D(\U4/Z_9 ), .CLK(clk), .Q(n14161), .QN(n12835) );
  DFFX1 \current_fsm_reg[10]  ( .D(\U4/Z_10 ), .CLK(clk), .QN(n11451) );
  DFFX1 \current_fsm_reg[11]  ( .D(\U4/Z_11 ), .CLK(clk), .QN(n11929) );
  DFFX1 \current_fsm_reg[12]  ( .D(\U4/Z_12 ), .CLK(clk), .QN(n12834) );
  DFFX1 \current_fsm_reg[13]  ( .D(\U4/Z_13 ), .CLK(clk), .QN(n11452) );
  DFFX1 \current_fsm_reg[14]  ( .D(\U4/Z_14 ), .CLK(clk), .QN(n11930) );
  DFFX1 \current_fsm_reg[15]  ( .D(\U4/Z_15 ), .CLK(clk), .Q(n13698), .QN(
        n12833) );
  DFFX1 \current_fsm_reg[16]  ( .D(\U4/Z_16 ), .CLK(clk), .QN(n11453) );
  DFFX1 \current_fsm_reg[17]  ( .D(\U4/Z_17 ), .CLK(clk), .QN(n11931) );
  DFFX1 \current_fsm_reg[18]  ( .D(\U4/Z_18 ), .CLK(clk), .QN(n12832) );
  DFFX1 \current_fsm_reg[19]  ( .D(\U4/Z_19 ), .CLK(clk), .QN(n11454) );
  DFFX1 \current_fsm_reg[20]  ( .D(\U4/Z_20 ), .CLK(clk), .QN(n11932) );
  DFFX1 \current_fsm_reg[21]  ( .D(\U4/Z_21 ), .CLK(clk), .Q(n14186), .QN(
        n11927) );
  DFFX1 \current_fsm_reg[22]  ( .D(\U4/Z_22 ), .CLK(clk), .QN(n11455) );
  DFFX1 \current_fsm_reg[23]  ( .D(\U4/Z_23 ), .CLK(clk), .QN(n11933) );
  DFFX1 \current_fsm_reg[24]  ( .D(\U4/Z_24 ), .CLK(clk), .QN(n12831) );
  DFFX1 \current_fsm_reg[25]  ( .D(\U4/Z_25 ), .CLK(clk), .QN(n11456) );
  DFFX1 \current_fsm_reg[26]  ( .D(\U4/Z_26 ), .CLK(clk), .QN(n11934) );
  DFFX1 \current_fsm_reg[27]  ( .D(\U4/Z_27 ), .CLK(clk), .QN(n12830) );
  DFFX1 \current_fsm_reg[28]  ( .D(\U4/Z_28 ), .CLK(clk), .QN(n11457) );
  DFFX1 \current_fsm_reg[29]  ( .D(\U4/Z_29 ), .CLK(clk), .Q(n11936) );
  DFFX1 \current_fsm_reg[30]  ( .D(\U4/Z_30 ), .CLK(clk), .Q(n13736), .QN(
        n11928) );
  DFFX1 \current_fsm_reg[31]  ( .D(\U4/Z_31 ), .CLK(clk), .QN(n11458) );
  DFFX1 \current_fsm_reg[32]  ( .D(\U4/Z_32 ), .CLK(clk), .Q(n11935) );
  DFFX1 \current_fsm_reg[33]  ( .D(\U4/Z_33 ), .CLK(clk), .QN(n11459) );
  DFFX1 \current_fsm_reg[34]  ( .D(\U4/Z_34 ), .CLK(clk), .QN(n11460) );
  DFFX1 \current_fsm_reg[35]  ( .D(\U4/Z_35 ), .CLK(clk), .Q(n14216), .QN(
        n12364) );
  DFFX1 \current_fsm_reg[36]  ( .D(\U4/Z_36 ), .CLK(clk), .Q(n14183), .QN(
        n12829) );
  DFFX1 \current_fsm_reg[37]  ( .D(\U4/Z_37 ), .CLK(clk), .QN(n11461) );
  DFFX1 \current_fsm_reg[38]  ( .D(\U4/Z_38 ), .CLK(clk), .QN(n11462) );
  DFFX1 \current_fsm_reg[39]  ( .D(\U4/Z_39 ), .CLK(clk), .Q(n14217), .QN(
        n12356) );
  DFFX1 \current_fsm_reg[41]  ( .D(\U4/Z_41 ), .CLK(clk), .QN(n11463) );
  DFFX1 \current_fsm_reg[42]  ( .D(\U4/Z_42 ), .CLK(clk), .QN(n11464) );
  DFFX1 \current_fsm_reg[44]  ( .D(\U4/Z_44 ), .CLK(clk), .QN(n11465) );
  DFFX1 \current_fsm_reg[45]  ( .D(\U4/Z_45 ), .CLK(clk), .QN(n12826) );
  DFFX1 \current_fsm_reg[47]  ( .D(\U4/Z_47 ), .CLK(clk), .QN(n11466) );
  DFFX1 \current_fsm_reg[51]  ( .D(\U4/Z_51 ), .CLK(clk), .QN(n11467) );
  DFFX1 \current_fsm_reg[52]  ( .D(\U4/Z_52 ), .CLK(clk), .QN(n11468) );
  DFFX1 \current_fsm_reg[54]  ( .D(\U4/Z_54 ), .CLK(clk), .QN(n11609) );
  DFFX1 \fmul_0_0_0_0_10_y_reg[11]  ( .D(n13137), .CLK(clk), .Q(n13916), .QN(
        n11655) );
  DFFX1 \fmul_0_0_0_0_10_y_reg[10]  ( .D(n13138), .CLK(clk), .Q(n13607), .QN(
        n11654) );
  DFFX1 \fmul_0_0_0_0_10_y_reg[9]  ( .D(n13139), .CLK(clk), .Q(n13967), .QN(
        n11653) );
  DFFX1 \fmul_0_0_0_0_10_y_reg[8]  ( .D(n13140), .CLK(clk), .Q(
        \fmul_0_0_0_0_10/add_2_root_add_321/B[4] ) );
  DFFX1 \fmul_0_0_0_0_10_y_reg[7]  ( .D(n13141), .CLK(clk), .Q(
        \fmul_0_0_0_0_10/add_2_root_add_321/B[3] ) );
  DFFX1 \fmul_0_0_0_0_10_y_reg[6]  ( .D(n13142), .CLK(clk), .Q(
        \fmul_0_0_0_0_10/add_2_root_add_321/B[2] ) );
  DFFX1 \fmul_0_0_0_0_10_y_reg[5]  ( .D(n13143), .CLK(clk), .Q(
        \fmul_0_0_0_0_10/add_2_root_add_321/B[1] ) );
  DFFX1 \fmul_0_0_0_0_10_y_reg[4]  ( .D(n13144), .CLK(clk), .Q(
        \fmul_0_0_0_0_10/add_2_root_add_321/B[0] ) );
  DFFX1 \fmul_0_0_0_0_10_y_reg[3]  ( .D(n13145), .CLK(clk), .Q(n13499), .QN(
        n12823) );
  DFFX1 \fmul_0_0_0_0_10_y_reg[2]  ( .D(n13146), .CLK(clk), .Q(n13617), .QN(
        n12824) );
  DFFX1 \fmul_0_0_0_0_10_y_reg[1]  ( .D(n13147), .CLK(clk), .Q(n13620), .QN(
        n12825) );
  DFFX1 \fmul_0_0_0_0_10_y_reg[0]  ( .D(n13148), .CLK(clk), .Q(n13618), .QN(
        n11923) );
  DFFX1 \fmul_0_0_0_0_9_y_reg[11]  ( .D(n13161), .CLK(clk), .Q(n13907), .QN(
        n11651) );
  DFFX1 \fmul_0_0_0_0_9_y_reg[10]  ( .D(n13162), .CLK(clk), .Q(n13606), .QN(
        n11650) );
  DFFX1 \fmul_0_0_0_0_9_y_reg[9]  ( .D(n13163), .CLK(clk), .Q(n13966), .QN(
        n11649) );
  DFFX1 \fmul_0_0_0_0_9_y_reg[8]  ( .D(n13164), .CLK(clk), .Q(n5302) );
  DFFX1 \fmul_0_0_0_0_9_y_reg[7]  ( .D(n13165), .CLK(clk), .Q(n5301) );
  DFFX1 \fmul_0_0_0_0_9_y_reg[6]  ( .D(n13166), .CLK(clk), .Q(n5300) );
  DFFX1 \fmul_0_0_0_0_9_y_reg[5]  ( .D(n13167), .CLK(clk), .Q(n5299) );
  DFFX1 \fmul_0_0_0_0_9_y_reg[4]  ( .D(n13168), .CLK(clk), .Q(n5298) );
  DFFX1 \fmul_0_0_0_0_9_y_reg[3]  ( .D(n13169), .CLK(clk), .Q(n5297) );
  DFFX1 \fmul_0_0_0_0_9_y_reg[2]  ( .D(n13170), .CLK(clk), .Q(n5296) );
  DFFX1 \fmul_0_0_0_0_9_y_reg[1]  ( .D(n13171), .CLK(clk), .Q(n5295) );
  DFFX1 \fmul_0_0_0_0_9_y_reg[0]  ( .D(n13172), .CLK(clk), .Q(n5294) );
  DFFX1 \fmul_0_0_0_0_8_y_reg[11]  ( .D(n13185), .CLK(clk), .Q(n13906), .QN(
        n11647) );
  DFFX1 \fmul_0_0_0_0_8_y_reg[10]  ( .D(n13186), .CLK(clk), .Q(n13605), .QN(
        n11646) );
  DFFX1 \fmul_0_0_0_0_8_y_reg[9]  ( .D(n13187), .CLK(clk), .Q(n13965), .QN(
        n11645) );
  DFFX1 \fmul_0_0_0_0_8_y_reg[8]  ( .D(n13188), .CLK(clk), .Q(n5374) );
  DFFX1 \fmul_0_0_0_0_8_y_reg[7]  ( .D(n13189), .CLK(clk), .Q(n5373) );
  DFFX1 \fmul_0_0_0_0_8_y_reg[6]  ( .D(n13190), .CLK(clk), .Q(n5372) );
  DFFX1 \fmul_0_0_0_0_8_y_reg[5]  ( .D(n13191), .CLK(clk), .Q(n5371) );
  DFFX1 \fmul_0_0_0_0_8_y_reg[4]  ( .D(n13192), .CLK(clk), .Q(n5370) );
  DFFX1 \fmul_0_0_0_0_8_y_reg[3]  ( .D(n13193), .CLK(clk), .Q(n5369) );
  DFFX1 \fmul_0_0_0_0_8_y_reg[2]  ( .D(n13194), .CLK(clk), .Q(n5368) );
  DFFX1 \fmul_0_0_0_0_8_y_reg[1]  ( .D(n13195), .CLK(clk), .Q(n5367) );
  DFFX1 \fmul_0_0_0_0_8_y_reg[0]  ( .D(n13196), .CLK(clk), .Q(n5366) );
  DFFX1 \fmul_0_0_0_0_7_y_reg[11]  ( .D(n13209), .CLK(clk), .Q(n13915), .QN(
        n11643) );
  DFFX1 \fmul_0_0_0_0_7_y_reg[10]  ( .D(n13210), .CLK(clk), .Q(n13905), .QN(
        n11642) );
  DFFX1 \fmul_0_0_0_0_7_y_reg[9]  ( .D(n13211), .CLK(clk), .Q(n14047), .QN(
        n11641) );
  DFFX1 \fmul_0_0_0_0_7_y_reg[8]  ( .D(n13212), .CLK(clk), .Q(n5446) );
  DFFX1 \fmul_0_0_0_0_7_y_reg[7]  ( .D(n13213), .CLK(clk), .Q(n5445) );
  DFFX1 \fmul_0_0_0_0_7_y_reg[6]  ( .D(n13214), .CLK(clk), .Q(n5444) );
  DFFX1 \fmul_0_0_0_0_7_y_reg[5]  ( .D(n13215), .CLK(clk), .Q(n5443) );
  DFFX1 \fmul_0_0_0_0_7_y_reg[4]  ( .D(n13216), .CLK(clk), .Q(n5442) );
  DFFX1 \fmul_0_0_0_0_7_y_reg[3]  ( .D(n13217), .CLK(clk), .Q(n5441) );
  DFFX1 \fmul_0_0_0_0_7_y_reg[2]  ( .D(n13218), .CLK(clk), .Q(n5440) );
  DFFX1 \fmul_0_0_0_0_7_y_reg[1]  ( .D(n13219), .CLK(clk), .Q(n5439) );
  DFFX1 \fmul_0_0_0_0_7_y_reg[0]  ( .D(n13220), .CLK(clk), .Q(n5438) );
  DFFX1 \fmul_0_0_0_0_6_y_reg[11]  ( .D(n13233), .CLK(clk), .Q(n13914), .QN(
        n11639) );
  DFFX1 \fmul_0_0_0_0_6_y_reg[10]  ( .D(n13234), .CLK(clk), .Q(n13904), .QN(
        n11638) );
  DFFX1 \fmul_0_0_0_0_6_y_reg[9]  ( .D(n13235), .CLK(clk), .Q(n14046), .QN(
        n11637) );
  DFFX1 \fmul_0_0_0_0_6_y_reg[8]  ( .D(n13236), .CLK(clk), .Q(n5518) );
  DFFX1 \fmul_0_0_0_0_6_y_reg[7]  ( .D(n13237), .CLK(clk), .Q(n5517) );
  DFFX1 \fmul_0_0_0_0_6_y_reg[6]  ( .D(n13238), .CLK(clk), .Q(n5516) );
  DFFX1 \fmul_0_0_0_0_6_y_reg[5]  ( .D(n13239), .CLK(clk), .Q(n5515) );
  DFFX1 \fmul_0_0_0_0_6_y_reg[4]  ( .D(n13240), .CLK(clk), .Q(n5514) );
  DFFX1 \fmul_0_0_0_0_6_y_reg[3]  ( .D(n13241), .CLK(clk), .Q(n5513) );
  DFFX1 \fmul_0_0_0_0_6_y_reg[2]  ( .D(n13242), .CLK(clk), .Q(n5512) );
  DFFX1 \fmul_0_0_0_0_6_y_reg[1]  ( .D(n13243), .CLK(clk), .Q(n5511) );
  DFFX1 \fmul_0_0_0_0_6_y_reg[0]  ( .D(n13244), .CLK(clk), .Q(n5510) );
  DFFX1 \fmul_0_0_0_0_5_y_reg[11]  ( .D(n13257), .CLK(clk), .Q(n13913), .QN(
        n11635) );
  DFFX1 \fmul_0_0_0_0_5_y_reg[10]  ( .D(n13258), .CLK(clk), .Q(n13903), .QN(
        n11634) );
  DFFX1 \fmul_0_0_0_0_5_y_reg[9]  ( .D(n13259), .CLK(clk), .Q(n14045), .QN(
        n11633) );
  DFFX1 \fmul_0_0_0_0_5_y_reg[8]  ( .D(n13260), .CLK(clk), .Q(n5590) );
  DFFX1 \fmul_0_0_0_0_5_y_reg[7]  ( .D(n13261), .CLK(clk), .Q(n5589) );
  DFFX1 \fmul_0_0_0_0_5_y_reg[6]  ( .D(n13262), .CLK(clk), .Q(n5588) );
  DFFX1 \fmul_0_0_0_0_5_y_reg[5]  ( .D(n13263), .CLK(clk), .Q(n5587) );
  DFFX1 \fmul_0_0_0_0_5_y_reg[4]  ( .D(n13264), .CLK(clk), .Q(n5586) );
  DFFX1 \fmul_0_0_0_0_5_y_reg[3]  ( .D(n13265), .CLK(clk), .Q(n5585) );
  DFFX1 \fmul_0_0_0_0_5_y_reg[2]  ( .D(n13266), .CLK(clk), .Q(n5584) );
  DFFX1 \fmul_0_0_0_0_5_y_reg[1]  ( .D(n13267), .CLK(clk), .Q(n5583) );
  DFFX1 \fmul_0_0_0_0_5_y_reg[0]  ( .D(n13268), .CLK(clk), .Q(n5582) );
  DFFX1 \fmul_0_0_0_0_4_y_reg[11]  ( .D(n13281), .CLK(clk), .Q(n13912), .QN(
        n11631) );
  DFFX1 \fmul_0_0_0_0_4_y_reg[10]  ( .D(n13282), .CLK(clk), .Q(n13902), .QN(
        n11630) );
  DFFX1 \fmul_0_0_0_0_4_y_reg[9]  ( .D(n13283), .CLK(clk), .Q(n14044), .QN(
        n11629) );
  DFFX1 \fmul_0_0_0_0_4_y_reg[8]  ( .D(n13284), .CLK(clk), .Q(n5662) );
  DFFX1 \fmul_0_0_0_0_4_y_reg[7]  ( .D(n13285), .CLK(clk), .Q(n5661) );
  DFFX1 \fmul_0_0_0_0_4_y_reg[6]  ( .D(n13286), .CLK(clk), .Q(n5660) );
  DFFX1 \fmul_0_0_0_0_4_y_reg[5]  ( .D(n13287), .CLK(clk), .Q(n5659) );
  DFFX1 \fmul_0_0_0_0_4_y_reg[4]  ( .D(n13288), .CLK(clk), .Q(n5658) );
  DFFX1 \fmul_0_0_0_0_4_y_reg[3]  ( .D(n13289), .CLK(clk), .Q(n5657) );
  DFFX1 \fmul_0_0_0_0_4_y_reg[2]  ( .D(n13290), .CLK(clk), .Q(n5656) );
  DFFX1 \fmul_0_0_0_0_4_y_reg[1]  ( .D(n13291), .CLK(clk), .Q(n5655) );
  DFFX1 \fmul_0_0_0_0_4_y_reg[0]  ( .D(n13292), .CLK(clk), .Q(n5654) );
  DFFX1 \fmul_0_0_0_0_3_y_reg[11]  ( .D(n13305), .CLK(clk), .Q(n13911), .QN(
        n11627) );
  DFFX1 \fmul_0_0_0_0_3_y_reg[10]  ( .D(n13306), .CLK(clk), .Q(n13901), .QN(
        n11626) );
  DFFX1 \fmul_0_0_0_0_3_y_reg[9]  ( .D(n13307), .CLK(clk), .Q(n14043), .QN(
        n11625) );
  DFFX1 \fmul_0_0_0_0_3_y_reg[8]  ( .D(n13308), .CLK(clk), .Q(n5734) );
  DFFX1 \fmul_0_0_0_0_3_y_reg[7]  ( .D(n13309), .CLK(clk), .Q(n5733) );
  DFFX1 \fmul_0_0_0_0_3_y_reg[6]  ( .D(n13310), .CLK(clk), .Q(n5732) );
  DFFX1 \fmul_0_0_0_0_3_y_reg[5]  ( .D(n13311), .CLK(clk), .Q(n5731) );
  DFFX1 \fmul_0_0_0_0_3_y_reg[4]  ( .D(n13312), .CLK(clk), .Q(n5730) );
  DFFX1 \fmul_0_0_0_0_3_y_reg[3]  ( .D(n13313), .CLK(clk), .Q(n5729) );
  DFFX1 \fmul_0_0_0_0_3_y_reg[2]  ( .D(n13314), .CLK(clk), .Q(n5728) );
  DFFX1 \fmul_0_0_0_0_3_y_reg[1]  ( .D(n13315), .CLK(clk), .Q(n5727) );
  DFFX1 \fmul_0_0_0_0_3_y_reg[0]  ( .D(n13316), .CLK(clk), .Q(n5726) );
  DFFX1 \fmul_0_0_0_0_2_y_reg[11]  ( .D(n13329), .CLK(clk), .Q(n13910), .QN(
        n11623) );
  DFFX1 \fmul_0_0_0_0_2_y_reg[10]  ( .D(n13330), .CLK(clk), .Q(n13900), .QN(
        n11622) );
  DFFX1 \fmul_0_0_0_0_2_y_reg[9]  ( .D(n13331), .CLK(clk), .Q(n14042), .QN(
        n11621) );
  DFFX1 \fmul_0_0_0_0_2_y_reg[8]  ( .D(n13332), .CLK(clk), .Q(n5806) );
  DFFX1 \fmul_0_0_0_0_2_y_reg[7]  ( .D(n13333), .CLK(clk), .Q(n5805) );
  DFFX1 \fmul_0_0_0_0_2_y_reg[6]  ( .D(n13334), .CLK(clk), .Q(n5804) );
  DFFX1 \fmul_0_0_0_0_2_y_reg[5]  ( .D(n13335), .CLK(clk), .Q(n5803) );
  DFFX1 \fmul_0_0_0_0_2_y_reg[4]  ( .D(n13336), .CLK(clk), .Q(n5802) );
  DFFX1 \fmul_0_0_0_0_2_y_reg[3]  ( .D(n13337), .CLK(clk), .Q(n5801) );
  DFFX1 \fmul_0_0_0_0_2_y_reg[2]  ( .D(n13338), .CLK(clk), .Q(n5800) );
  DFFX1 \fmul_0_0_0_0_2_y_reg[1]  ( .D(n13339), .CLK(clk), .Q(n5799) );
  DFFX1 \fmul_0_0_0_0_2_y_reg[0]  ( .D(n13340), .CLK(clk), .Q(n5798) );
  DFFX1 \fmul_0_0_0_0_1_y_reg[11]  ( .D(n13353), .CLK(clk), .Q(n13909), .QN(
        n11619) );
  DFFX1 \fmul_0_0_0_0_1_y_reg[10]  ( .D(n13354), .CLK(clk), .Q(n13899), .QN(
        n11618) );
  DFFX1 \fmul_0_0_0_0_1_y_reg[9]  ( .D(n13355), .CLK(clk), .Q(n14041), .QN(
        n11617) );
  DFFX1 \fmul_0_0_0_0_1_y_reg[8]  ( .D(n13356), .CLK(clk), .Q(n5878) );
  DFFX1 \fmul_0_0_0_0_1_y_reg[7]  ( .D(n13357), .CLK(clk), .Q(n5877) );
  DFFX1 \fmul_0_0_0_0_1_y_reg[6]  ( .D(n13358), .CLK(clk), .Q(n5876) );
  DFFX1 \fmul_0_0_0_0_1_y_reg[5]  ( .D(n13359), .CLK(clk), .Q(n5875) );
  DFFX1 \fmul_0_0_0_0_1_y_reg[4]  ( .D(n13360), .CLK(clk), .Q(n5874) );
  DFFX1 \fmul_0_0_0_0_1_y_reg[3]  ( .D(n13361), .CLK(clk), .Q(n5873) );
  DFFX1 \fmul_0_0_0_0_1_y_reg[2]  ( .D(n13362), .CLK(clk), .Q(n5872) );
  DFFX1 \fmul_0_0_0_0_1_y_reg[1]  ( .D(n13363), .CLK(clk), .Q(n5871) );
  DFFX1 \fmul_0_0_0_0_1_y_reg[0]  ( .D(n13364), .CLK(clk), .Q(n5870) );
  DFFX1 \fmul_0_0_0_0_0_y_reg[11]  ( .D(n13376), .CLK(clk), .Q(n13908), .QN(
        n11615) );
  DFFX1 \fmul_0_0_0_0_0_y_reg[10]  ( .D(n13377), .CLK(clk), .Q(n13898), .QN(
        n11614) );
  DFFX1 \fmul_0_0_0_0_0_y_reg[9]  ( .D(n13378), .CLK(clk), .Q(n14040), .QN(
        n11613) );
  DFFX1 \fmul_0_0_0_0_0_y_reg[8]  ( .D(n13379), .CLK(clk), .Q(n5950) );
  DFFX1 \fmul_0_0_0_0_0_y_reg[7]  ( .D(n13380), .CLK(clk), .Q(n5949) );
  DFFX1 \fmul_0_0_0_0_0_y_reg[6]  ( .D(n13381), .CLK(clk), .Q(n5948) );
  DFFX1 \fmul_0_0_0_0_0_y_reg[5]  ( .D(n13382), .CLK(clk), .Q(n5947) );
  DFFX1 \fmul_0_0_0_0_0_y_reg[4]  ( .D(n13383), .CLK(clk), .Q(n5946) );
  DFFX1 \fmul_0_0_0_0_0_y_reg[3]  ( .D(n13384), .CLK(clk), .Q(n5945) );
  DFFX1 \fmul_0_0_0_0_0_y_reg[2]  ( .D(n13385), .CLK(clk), .Q(n5944) );
  DFFX1 \fmul_0_0_0_0_0_y_reg[1]  ( .D(n13386), .CLK(clk), .Q(n5943) );
  DFFX1 \fmul_0_0_0_0_0_y_reg[0]  ( .D(n13387), .CLK(clk), .Q(n5942) );
  DFFX1 \fmul_0_0_0_0_10_x_reg[11]  ( .D(n13149), .CLK(clk), .Q(n13765), .QN(
        n12815) );
  DFFX1 \fmul_0_0_0_0_9_x_reg[11]  ( .D(n13173), .CLK(clk), .Q(n13764), .QN(
        n12787) );
  DFFX1 \fmul_0_0_0_0_8_x_reg[11]  ( .D(n13197), .CLK(clk), .Q(n13763), .QN(
        n12777) );
  DFFX1 \fmul_0_0_0_0_7_x_reg[11]  ( .D(n13221), .CLK(clk), .Q(n13762), .QN(
        n12767) );
  DFFX1 \fmul_0_0_0_0_6_x_reg[11]  ( .D(n13245), .CLK(clk), .Q(n13761), .QN(
        n12749) );
  DFFX1 \fmul_0_0_0_0_5_x_reg[11]  ( .D(n13269), .CLK(clk), .Q(n13760), .QN(
        n12747) );
  DFFX1 \fmul_0_0_0_0_4_x_reg[11]  ( .D(n13293), .CLK(clk), .Q(n13759), .QN(
        n12729) );
  DFFX1 \fmul_0_0_0_0_3_x_reg[11]  ( .D(n13317), .CLK(clk), .Q(n13758), .QN(
        n12727) );
  DFFX1 \fmul_0_0_0_0_2_x_reg[11]  ( .D(n13341), .CLK(clk), .Q(n13757), .QN(
        n12709) );
  DFFX1 \fmul_0_0_0_0_1_x_reg[11]  ( .D(n13365), .CLK(clk), .Q(n13756), .QN(
        n12707) );
  DFFX1 \fmul_0_0_0_0_0_x_reg[11]  ( .D(n13388), .CLK(clk), .Q(n13755), .QN(
        n12689) );
  DFFX1 \fmul_0_0_0_0_10_x_reg[10]  ( .D(n13150), .CLK(clk), .Q(n13897), .QN(
        n12816) );
  DFFX1 \fmul_0_0_0_0_9_x_reg[10]  ( .D(n13174), .CLK(clk), .Q(n13896), .QN(
        n12788) );
  DFFX1 \fmul_0_0_0_0_8_x_reg[10]  ( .D(n13198), .CLK(clk), .Q(n13895), .QN(
        n12778) );
  DFFX1 \fmul_0_0_0_0_7_x_reg[10]  ( .D(n13222), .CLK(clk), .Q(n13615), .QN(
        n12768) );
  DFFX1 \fmul_0_0_0_0_6_x_reg[10]  ( .D(n13246), .CLK(clk), .Q(n13614), .QN(
        n12750) );
  DFFX1 \fmul_0_0_0_0_5_x_reg[10]  ( .D(n13270), .CLK(clk), .Q(n13613), .QN(
        n12748) );
  DFFX1 \fmul_0_0_0_0_4_x_reg[10]  ( .D(n13294), .CLK(clk), .Q(n13612), .QN(
        n12730) );
  DFFX1 \fmul_0_0_0_0_3_x_reg[10]  ( .D(n13318), .CLK(clk), .Q(n13611), .QN(
        n12728) );
  DFFX1 \fmul_0_0_0_0_2_x_reg[10]  ( .D(n13342), .CLK(clk), .Q(n13610), .QN(
        n12710) );
  DFFX1 \fmul_0_0_0_0_1_x_reg[10]  ( .D(n13366), .CLK(clk), .Q(n13609), .QN(
        n12708) );
  DFFX1 \fmul_0_0_0_0_0_x_reg[10]  ( .D(n13389), .CLK(clk), .Q(n13608), .QN(
        n12690) );
  DFFX1 \fmul_0_0_0_0_10_x_reg[9]  ( .D(n13151), .CLK(clk), .Q(n14077), .QN(
        n11652) );
  DFFX1 \fmul_0_0_0_0_9_x_reg[9]  ( .D(n13175), .CLK(clk), .Q(n14076), .QN(
        n11648) );
  DFFX1 \fmul_0_0_0_0_8_x_reg[9]  ( .D(n13199), .CLK(clk), .Q(n14075), .QN(
        n11644) );
  DFFX1 \fmul_0_0_0_0_7_x_reg[9]  ( .D(n13223), .CLK(clk), .Q(n14074), .QN(
        n11640) );
  DFFX1 \fmul_0_0_0_0_6_x_reg[9]  ( .D(n13247), .CLK(clk), .Q(n14073), .QN(
        n11636) );
  DFFX1 \fmul_0_0_0_0_5_x_reg[9]  ( .D(n13271), .CLK(clk), .Q(n14072), .QN(
        n11632) );
  DFFX1 \fmul_0_0_0_0_4_x_reg[9]  ( .D(n13295), .CLK(clk), .Q(n14071), .QN(
        n11628) );
  DFFX1 \fmul_0_0_0_0_3_x_reg[9]  ( .D(n13319), .CLK(clk), .Q(n14070), .QN(
        n11624) );
  DFFX1 \fmul_0_0_0_0_2_x_reg[9]  ( .D(n13343), .CLK(clk), .Q(n14069), .QN(
        n11620) );
  DFFX1 \fmul_0_0_0_0_1_x_reg[9]  ( .D(n13367), .CLK(clk), .Q(n14068), .QN(
        n11616) );
  DFFX1 \fmul_0_0_0_0_0_x_reg[9]  ( .D(n13390), .CLK(clk), .Q(n14067), .QN(
        n11612) );
  DFFX1 \fmul_0_0_0_0_10_x_reg[8]  ( .D(n13152), .CLK(clk), .Q(
        \fmul_0_0_0_0_10/add_2_root_add_321/A[4] ) );
  DFFX1 \fmul_0_0_0_0_9_x_reg[8]  ( .D(n13176), .CLK(clk), .Q(n5314) );
  DFFX1 \fmul_0_0_0_0_8_x_reg[8]  ( .D(n13200), .CLK(clk), .Q(n5386) );
  DFFX1 \fmul_0_0_0_0_7_x_reg[8]  ( .D(n13224), .CLK(clk), .Q(n5458) );
  DFFX1 \fmul_0_0_0_0_6_x_reg[8]  ( .D(n13248), .CLK(clk), .Q(n5530) );
  DFFX1 \fmul_0_0_0_0_5_x_reg[8]  ( .D(n13272), .CLK(clk), .Q(n5602) );
  DFFX1 \fmul_0_0_0_0_4_x_reg[8]  ( .D(n13296), .CLK(clk), .Q(n5674) );
  DFFX1 \fmul_0_0_0_0_3_x_reg[8]  ( .D(n13320), .CLK(clk), .Q(n5746) );
  DFFX1 \fmul_0_0_0_0_2_x_reg[8]  ( .D(n13344), .CLK(clk), .Q(n5818) );
  DFFX1 \fmul_0_0_0_0_1_x_reg[8]  ( .D(n13368), .CLK(clk), .Q(n5890) );
  DFFX1 \fmul_0_0_0_0_0_x_reg[8]  ( .D(n13391), .CLK(clk), .Q(n5962) );
  DFFX1 \fmul_0_0_0_0_10_x_reg[7]  ( .D(n13153), .CLK(clk), .Q(
        \fmul_0_0_0_0_10/add_2_root_add_321/A[3] ) );
  DFFX1 \fmul_0_0_0_0_9_x_reg[7]  ( .D(n13177), .CLK(clk), .Q(n5313) );
  DFFX1 \fmul_0_0_0_0_8_x_reg[7]  ( .D(n13201), .CLK(clk), .Q(n5385) );
  DFFX1 \fmul_0_0_0_0_7_x_reg[7]  ( .D(n13225), .CLK(clk), .Q(n5457) );
  DFFX1 \fmul_0_0_0_0_6_x_reg[7]  ( .D(n13249), .CLK(clk), .Q(n5529) );
  DFFX1 \fmul_0_0_0_0_5_x_reg[7]  ( .D(n13273), .CLK(clk), .Q(n5601) );
  DFFX1 \fmul_0_0_0_0_4_x_reg[7]  ( .D(n13297), .CLK(clk), .Q(n5673) );
  DFFX1 \fmul_0_0_0_0_3_x_reg[7]  ( .D(n13321), .CLK(clk), .Q(n5745) );
  DFFX1 \fmul_0_0_0_0_2_x_reg[7]  ( .D(n13345), .CLK(clk), .Q(n5817) );
  DFFX1 \fmul_0_0_0_0_1_x_reg[7]  ( .D(n13369), .CLK(clk), .Q(n5889) );
  DFFX1 \fmul_0_0_0_0_0_x_reg[7]  ( .D(n13392), .CLK(clk), .Q(n5961) );
  DFFX1 \fmul_0_0_0_0_10_x_reg[6]  ( .D(n13154), .CLK(clk), .Q(
        \fmul_0_0_0_0_10/add_2_root_add_321/A[2] ) );
  DFFX1 \fmul_0_0_0_0_9_x_reg[6]  ( .D(n13178), .CLK(clk), .Q(n5312) );
  DFFX1 \fmul_0_0_0_0_8_x_reg[6]  ( .D(n13202), .CLK(clk), .Q(n5384) );
  DFFX1 \fmul_0_0_0_0_7_x_reg[6]  ( .D(n13226), .CLK(clk), .Q(n5456) );
  DFFX1 \fmul_0_0_0_0_6_x_reg[6]  ( .D(n13250), .CLK(clk), .Q(n5528) );
  DFFX1 \fmul_0_0_0_0_5_x_reg[6]  ( .D(n13274), .CLK(clk), .Q(n5600) );
  DFFX1 \fmul_0_0_0_0_4_x_reg[6]  ( .D(n13298), .CLK(clk), .Q(n5672) );
  DFFX1 \fmul_0_0_0_0_3_x_reg[6]  ( .D(n13322), .CLK(clk), .Q(n5744) );
  DFFX1 \fmul_0_0_0_0_2_x_reg[6]  ( .D(n13346), .CLK(clk), .Q(n5816) );
  DFFX1 \fmul_0_0_0_0_1_x_reg[6]  ( .D(n13370), .CLK(clk), .Q(n5888) );
  DFFX1 \fmul_0_0_0_0_0_x_reg[6]  ( .D(n13393), .CLK(clk), .Q(n5960) );
  DFFX1 \fmul_0_0_0_0_10_x_reg[5]  ( .D(n13155), .CLK(clk), .Q(
        \fmul_0_0_0_0_10/add_2_root_add_321/A[1] ) );
  DFFX1 \fmul_0_0_0_0_9_x_reg[5]  ( .D(n13179), .CLK(clk), .Q(n5311) );
  DFFX1 \fmul_0_0_0_0_8_x_reg[5]  ( .D(n13203), .CLK(clk), .Q(n5383) );
  DFFX1 \fmul_0_0_0_0_7_x_reg[5]  ( .D(n13227), .CLK(clk), .Q(n5455) );
  DFFX1 \fmul_0_0_0_0_6_x_reg[5]  ( .D(n13251), .CLK(clk), .Q(n5527) );
  DFFX1 \fmul_0_0_0_0_5_x_reg[5]  ( .D(n13275), .CLK(clk), .Q(n5599) );
  DFFX1 \fmul_0_0_0_0_4_x_reg[5]  ( .D(n13299), .CLK(clk), .Q(n5671) );
  DFFX1 \fmul_0_0_0_0_3_x_reg[5]  ( .D(n13323), .CLK(clk), .Q(n5743) );
  DFFX1 \fmul_0_0_0_0_2_x_reg[5]  ( .D(n13347), .CLK(clk), .Q(n5815) );
  DFFX1 \fmul_0_0_0_0_1_x_reg[5]  ( .D(n13371), .CLK(clk), .Q(n5887) );
  DFFX1 \fmul_0_0_0_0_0_x_reg[5]  ( .D(n13394), .CLK(clk), .Q(n5959) );
  DFFX1 \fmul_0_0_0_0_10_x_reg[4]  ( .D(n13156), .CLK(clk), .Q(
        \fmul_0_0_0_0_10/add_2_root_add_321/A[0] ) );
  DFFX1 \fmul_0_0_0_0_9_x_reg[4]  ( .D(n13180), .CLK(clk), .Q(n5310) );
  DFFX1 \fmul_0_0_0_0_8_x_reg[4]  ( .D(n13204), .CLK(clk), .Q(n5382) );
  DFFX1 \fmul_0_0_0_0_7_x_reg[4]  ( .D(n13228), .CLK(clk), .Q(n5454) );
  DFFX1 \fmul_0_0_0_0_6_x_reg[4]  ( .D(n13252), .CLK(clk), .Q(n5526) );
  DFFX1 \fmul_0_0_0_0_5_x_reg[4]  ( .D(n13276), .CLK(clk), .Q(n5598) );
  DFFX1 \fmul_0_0_0_0_4_x_reg[4]  ( .D(n13300), .CLK(clk), .Q(n5670) );
  DFFX1 \fmul_0_0_0_0_3_x_reg[4]  ( .D(n13324), .CLK(clk), .Q(n5742) );
  DFFX1 \fmul_0_0_0_0_2_x_reg[4]  ( .D(n13348), .CLK(clk), .Q(n5814) );
  DFFX1 \fmul_0_0_0_0_1_x_reg[4]  ( .D(n13372), .CLK(clk), .Q(n5886) );
  DFFX1 \fmul_0_0_0_0_0_x_reg[4]  ( .D(n13395), .CLK(clk), .Q(n5958) );
  DFFX1 \fmul_0_0_0_0_10_x_reg[3]  ( .D(n13157), .CLK(clk), .Q(n13468), .QN(
        n11924) );
  DFFX1 \fmul_0_0_0_0_9_x_reg[3]  ( .D(n13181), .CLK(clk), .Q(n5309) );
  DFFX1 \fmul_0_0_0_0_8_x_reg[3]  ( .D(n13205), .CLK(clk), .Q(n5381) );
  DFFX1 \fmul_0_0_0_0_7_x_reg[3]  ( .D(n13229), .CLK(clk), .Q(n5453) );
  DFFX1 \fmul_0_0_0_0_6_x_reg[3]  ( .D(n13253), .CLK(clk), .Q(n5525) );
  DFFX1 \fmul_0_0_0_0_5_x_reg[3]  ( .D(n13277), .CLK(clk), .Q(n5597) );
  DFFX1 \fmul_0_0_0_0_4_x_reg[3]  ( .D(n13301), .CLK(clk), .Q(n5669) );
  DFFX1 \fmul_0_0_0_0_3_x_reg[3]  ( .D(n13325), .CLK(clk), .Q(n5741) );
  DFFX1 \fmul_0_0_0_0_2_x_reg[3]  ( .D(n13349), .CLK(clk), .Q(n5813) );
  DFFX1 \fmul_0_0_0_0_1_x_reg[3]  ( .D(n13373), .CLK(clk), .Q(n5885) );
  DFFX1 \fmul_0_0_0_0_0_x_reg[3]  ( .D(n13396), .CLK(clk), .Q(n5957) );
  DFFX1 \fmul_0_0_0_0_10_x_reg[2]  ( .D(n13158), .CLK(clk), .Q(n13619), .QN(
        n12820) );
  DFFX1 \fmul_0_0_0_0_9_x_reg[2]  ( .D(n13182), .CLK(clk), .Q(n5308) );
  DFFX1 \fmul_0_0_0_0_8_x_reg[2]  ( .D(n13206), .CLK(clk), .Q(n5380) );
  DFFX1 \fmul_0_0_0_0_7_x_reg[2]  ( .D(n13230), .CLK(clk), .Q(n5452) );
  DFFX1 \fmul_0_0_0_0_6_x_reg[2]  ( .D(n13254), .CLK(clk), .Q(n5524) );
  DFFX1 \fmul_0_0_0_0_5_x_reg[2]  ( .D(n13278), .CLK(clk), .Q(n5596) );
  DFFX1 \fmul_0_0_0_0_4_x_reg[2]  ( .D(n13302), .CLK(clk), .Q(n5668) );
  DFFX1 \fmul_0_0_0_0_3_x_reg[2]  ( .D(n13326), .CLK(clk), .Q(n5740) );
  DFFX1 \fmul_0_0_0_0_2_x_reg[2]  ( .D(n13350), .CLK(clk), .Q(n5812) );
  DFFX1 \fmul_0_0_0_0_1_x_reg[2]  ( .D(n13374), .CLK(clk), .Q(n5884) );
  DFFX1 \fmul_0_0_0_0_0_x_reg[2]  ( .D(n13397), .CLK(clk), .Q(n5956) );
  DFFX1 \fmul_0_0_0_0_10_x_reg[1]  ( .D(n13159), .CLK(clk), .Q(n13629), .QN(
        n12821) );
  DFFX1 \fmul_0_0_0_0_9_x_reg[1]  ( .D(n13183), .CLK(clk), .Q(n5307) );
  DFFX1 \fmul_0_0_0_0_8_x_reg[1]  ( .D(n13207), .CLK(clk), .Q(n5379) );
  DFFX1 \fmul_0_0_0_0_7_x_reg[1]  ( .D(n13231), .CLK(clk), .Q(n5451) );
  DFFX1 \fmul_0_0_0_0_6_x_reg[1]  ( .D(n13255), .CLK(clk), .Q(n5523) );
  DFFX1 \fmul_0_0_0_0_5_x_reg[1]  ( .D(n13279), .CLK(clk), .Q(n5595) );
  DFFX1 \fmul_0_0_0_0_4_x_reg[1]  ( .D(n13303), .CLK(clk), .Q(n5667) );
  DFFX1 \fmul_0_0_0_0_3_x_reg[1]  ( .D(n13327), .CLK(clk), .Q(n5739) );
  DFFX1 \fmul_0_0_0_0_2_x_reg[1]  ( .D(n13351), .CLK(clk), .Q(n5811) );
  DFFX1 \fmul_0_0_0_0_1_x_reg[1]  ( .D(n13375), .CLK(clk), .Q(n5883) );
  DFFX1 \fmul_0_0_0_0_0_x_reg[1]  ( .D(n13398), .CLK(clk), .Q(n5955) );
  DFFX1 \fmul_0_0_0_0_10_x_reg[0]  ( .D(n13136), .CLK(clk), .Q(n13498), .QN(
        n12822) );
  DFFX1 \fmul_0_0_0_0_9_x_reg[0]  ( .D(n13160), .CLK(clk), .Q(n5306) );
  DFFX1 \fmul_0_0_0_0_8_x_reg[0]  ( .D(n13184), .CLK(clk), .Q(n5378) );
  DFFX1 \fmul_0_0_0_0_7_x_reg[0]  ( .D(n13208), .CLK(clk), .Q(n5450) );
  DFFX1 \fmul_0_0_0_0_6_x_reg[0]  ( .D(n13232), .CLK(clk), .Q(n5522) );
  DFFX1 \fmul_0_0_0_0_5_x_reg[0]  ( .D(n13256), .CLK(clk), .Q(n5594) );
  DFFX1 \fmul_0_0_0_0_4_x_reg[0]  ( .D(n13280), .CLK(clk), .Q(n5666) );
  DFFX1 \fmul_0_0_0_0_3_x_reg[0]  ( .D(n13304), .CLK(clk), .Q(n5738) );
  DFFX1 \fmul_0_0_0_0_2_x_reg[0]  ( .D(n13328), .CLK(clk), .Q(n5810) );
  DFFX1 \fmul_0_0_0_0_1_x_reg[0]  ( .D(n13352), .CLK(clk), .Q(n5882) );
  DFFX1 \fmul_0_0_0_0_0_x_reg[0]  ( .D(n13399), .CLK(clk), .Q(n5954) );
  DFFX1 \fadd_0_0_0_0_0/norm/n351_q_reg[0]  ( .D(
        \fadd_0_0_0_0_0/fracrclose1 [0]), .CLK(clk), .QN(n11471) );
  DFFX1 \fadd_0_0_0_0_0/norm/n351_q_reg[1]  ( .D(
        \fadd_0_0_0_0_0/fracrclose1 [1]), .CLK(clk), .QN(n11472) );
  DFFX1 \fadd_0_0_0_0_0/norm/n351_q_reg[2]  ( .D(
        \fadd_0_0_0_0_0/fracrclose1 [2]), .CLK(clk), .Q(n14048), .QN(n11882)
         );
  DFFX1 \fadd_0_0_0_0_0/norm/n351_q_reg[3]  ( .D(
        \fadd_0_0_0_0_0/fracrclose1 [3]), .CLK(clk), .QN(n11881) );
  DFFX1 \fadd_0_0_0_0_0/norm/n351_q_reg[4]  ( .D(
        \fadd_0_0_0_0_0/fracrclose1 [4]), .CLK(clk), .QN(n11880) );
  DFFX1 \fadd_0_0_0_0_0/norm/n351_q_reg[5]  ( .D(
        \fadd_0_0_0_0_0/fracrclose1 [5]), .CLK(clk), .Q(n13548), .QN(n11879)
         );
  DFFX1 \fadd_0_0_0_0_0/norm/n352_q_reg[4]  ( .D(
        \fadd_0_0_0_0_0/norm/level1 [4]), .CLK(clk), .Q(
        \fadd_0_0_0_0_0/norm/level1_d1[4] ) );
  DFFX1 \fadd_0_0_0_0_0/norm/n353_q_reg  ( .D(\fadd_0_0_0_0_0/sub_784/B[0] ), 
        .CLK(clk), .QN(n12849) );
  DFFX1 \fadd_0_0_0_0_0/norm/n352_q_reg[3]  ( .D(
        \fadd_0_0_0_0_0/norm/level1 [3]), .CLK(clk), .Q(n13700) );
  DFFX1 \fadd_0_0_0_0_0/norm/n352_q_reg[2]  ( .D(
        \fadd_0_0_0_0_0/norm/level1 [2]), .CLK(clk), .Q(n13564) );
  DFFX1 \fadd_0_0_0_0_0/norm/n352_q_reg[1]  ( .D(
        \fadd_0_0_0_0_0/norm/level1 [1]), .CLK(clk), .Q(n13487) );
  DFFX1 \fadd_0_0_0_0_0/norm/n352_q_reg[0]  ( .D(
        \fadd_0_0_0_0_0/norm/level1 [0]), .CLK(clk), .Q(n13679) );
  DFFX1 \fadd_0_0_0_0_1/norm/n351_q_reg[0]  ( .D(
        \fadd_0_0_0_0_1/fracrclose1 [0]), .CLK(clk), .QN(n11484) );
  DFFX1 \fadd_0_0_0_0_1/norm/n351_q_reg[1]  ( .D(
        \fadd_0_0_0_0_1/fracrclose1 [1]), .CLK(clk), .QN(n11485) );
  DFFX1 \fadd_0_0_0_0_1/norm/n351_q_reg[2]  ( .D(
        \fadd_0_0_0_0_1/fracrclose1 [2]), .CLK(clk), .Q(n14049), .QN(n11886)
         );
  DFFX1 \fadd_0_0_0_0_1/norm/n351_q_reg[3]  ( .D(
        \fadd_0_0_0_0_1/fracrclose1 [3]), .CLK(clk), .QN(n11885) );
  DFFX1 \fadd_0_0_0_0_1/norm/n351_q_reg[4]  ( .D(
        \fadd_0_0_0_0_1/fracrclose1 [4]), .CLK(clk), .QN(n11884) );
  DFFX1 \fadd_0_0_0_0_1/norm/n351_q_reg[5]  ( .D(
        \fadd_0_0_0_0_1/fracrclose1 [5]), .CLK(clk), .Q(n13547), .QN(n11883)
         );
  DFFX1 \fadd_0_0_0_0_1/norm/n352_q_reg[4]  ( .D(
        \fadd_0_0_0_0_1/norm/level1 [4]), .CLK(clk), .Q(
        \fadd_0_0_0_0_1/norm/level1_d1[4] ) );
  DFFX1 \fadd_0_0_0_0_1/norm/n353_q_reg  ( .D(\fadd_0_0_0_0_1/sub_784/B[0] ), 
        .CLK(clk), .QN(n12851) );
  DFFX1 \fadd_0_0_0_0_1/norm/n352_q_reg[3]  ( .D(
        \fadd_0_0_0_0_1/norm/level1 [3]), .CLK(clk), .Q(n13701) );
  DFFX1 \fadd_0_0_0_0_1/norm/n352_q_reg[2]  ( .D(
        \fadd_0_0_0_0_1/norm/level1 [2]), .CLK(clk), .Q(n13565) );
  DFFX1 \fadd_0_0_0_0_1/norm/n352_q_reg[1]  ( .D(
        \fadd_0_0_0_0_1/norm/level1 [1]), .CLK(clk), .Q(n13488) );
  DFFX1 \fadd_0_0_0_0_1/norm/n352_q_reg[0]  ( .D(
        \fadd_0_0_0_0_1/norm/level1 [0]), .CLK(clk), .Q(n13680) );
  DFFX1 \fadd_0_0_0_0_2/norm/n351_q_reg[0]  ( .D(
        \fadd_0_0_0_0_2/fracrclose1 [0]), .CLK(clk), .QN(n11506) );
  DFFX1 \fadd_0_0_0_0_2/norm/n351_q_reg[1]  ( .D(
        \fadd_0_0_0_0_2/fracrclose1 [1]), .CLK(clk), .QN(n11507) );
  DFFX1 \fadd_0_0_0_0_2/norm/n351_q_reg[2]  ( .D(
        \fadd_0_0_0_0_2/fracrclose1 [2]), .CLK(clk), .Q(n14050), .QN(n11894)
         );
  DFFX1 \fadd_0_0_0_0_2/norm/n351_q_reg[3]  ( .D(
        \fadd_0_0_0_0_2/fracrclose1 [3]), .CLK(clk), .QN(n11893) );
  DFFX1 \fadd_0_0_0_0_2/norm/n351_q_reg[4]  ( .D(
        \fadd_0_0_0_0_2/fracrclose1 [4]), .CLK(clk), .QN(n11892) );
  DFFX1 \fadd_0_0_0_0_2/norm/n351_q_reg[5]  ( .D(
        \fadd_0_0_0_0_2/fracrclose1 [5]), .CLK(clk), .Q(n13546), .QN(n11891)
         );
  DFFX1 \fadd_0_0_0_0_2/norm/n352_q_reg[4]  ( .D(
        \fadd_0_0_0_0_2/norm/level1 [4]), .CLK(clk), .Q(
        \fadd_0_0_0_0_2/norm/level1_d1[4] ) );
  DFFX1 \fadd_0_0_0_0_2/norm/n353_q_reg  ( .D(\fadd_0_0_0_0_2/sub_784/B[0] ), 
        .CLK(clk), .QN(n12853) );
  DFFX1 \fadd_0_0_0_0_2/norm/n352_q_reg[3]  ( .D(
        \fadd_0_0_0_0_2/norm/level1 [3]), .CLK(clk), .Q(n13694) );
  DFFX1 \fadd_0_0_0_0_2/norm/n352_q_reg[2]  ( .D(
        \fadd_0_0_0_0_2/norm/level1 [2]), .CLK(clk), .Q(n13552) );
  DFFX1 \fadd_0_0_0_0_2/norm/n352_q_reg[1]  ( .D(
        \fadd_0_0_0_0_2/norm/level1 [1]), .CLK(clk), .Q(n13484) );
  DFFX1 \fadd_0_0_0_0_2/norm/n352_q_reg[0]  ( .D(
        \fadd_0_0_0_0_2/norm/level1 [0]), .CLK(clk), .Q(n13675) );
  DFFX1 \fadd_0_0_0_0_3/norm/n351_q_reg[0]  ( .D(
        \fadd_0_0_0_0_3/fracrclose1 [0]), .CLK(clk), .QN(n11519) );
  DFFX1 \fadd_0_0_0_0_3/norm/n351_q_reg[1]  ( .D(
        \fadd_0_0_0_0_3/fracrclose1 [1]), .CLK(clk), .QN(n11520) );
  DFFX1 \fadd_0_0_0_0_3/norm/n351_q_reg[2]  ( .D(
        \fadd_0_0_0_0_3/fracrclose1 [2]), .CLK(clk), .Q(n14051), .QN(n11898)
         );
  DFFX1 \fadd_0_0_0_0_3/norm/n351_q_reg[3]  ( .D(
        \fadd_0_0_0_0_3/fracrclose1 [3]), .CLK(clk), .QN(n11897) );
  DFFX1 \fadd_0_0_0_0_3/norm/n351_q_reg[4]  ( .D(
        \fadd_0_0_0_0_3/fracrclose1 [4]), .CLK(clk), .QN(n11896) );
  DFFX1 \fadd_0_0_0_0_3/norm/n351_q_reg[5]  ( .D(
        \fadd_0_0_0_0_3/fracrclose1 [5]), .CLK(clk), .Q(n13545), .QN(n11895)
         );
  DFFX1 \fadd_0_0_0_0_3/norm/n352_q_reg[4]  ( .D(
        \fadd_0_0_0_0_3/norm/level1 [4]), .CLK(clk), .Q(
        \fadd_0_0_0_0_3/norm/level1_d1[4] ) );
  DFFX1 \fadd_0_0_0_0_3/norm/n353_q_reg  ( .D(\fadd_0_0_0_0_3/sub_784/B[0] ), 
        .CLK(clk), .QN(n12855) );
  DFFX1 \fadd_0_0_0_0_3/norm/n352_q_reg[3]  ( .D(
        \fadd_0_0_0_0_3/norm/level1 [3]), .CLK(clk), .Q(n13702) );
  DFFX1 \fadd_0_0_0_0_3/norm/n352_q_reg[2]  ( .D(
        \fadd_0_0_0_0_3/norm/level1 [2]), .CLK(clk), .Q(n13566) );
  DFFX1 \fadd_0_0_0_0_3/norm/n352_q_reg[1]  ( .D(
        \fadd_0_0_0_0_3/norm/level1 [1]), .CLK(clk), .Q(n13489) );
  DFFX1 \fadd_0_0_0_0_3/norm/n352_q_reg[0]  ( .D(
        \fadd_0_0_0_0_3/norm/level1 [0]), .CLK(clk), .Q(n13681) );
  DFFX1 \fadd_0_0_0_0_4/norm/n351_q_reg[0]  ( .D(
        \fadd_0_0_0_0_4/fracrclose1 [0]), .CLK(clk), .QN(n11532) );
  DFFX1 \fadd_0_0_0_0_4/norm/n351_q_reg[1]  ( .D(
        \fadd_0_0_0_0_4/fracrclose1 [1]), .CLK(clk), .QN(n11533) );
  DFFX1 \fadd_0_0_0_0_4/norm/n351_q_reg[2]  ( .D(
        \fadd_0_0_0_0_4/fracrclose1 [2]), .CLK(clk), .Q(n14052), .QN(n11902)
         );
  DFFX1 \fadd_0_0_0_0_4/norm/n351_q_reg[3]  ( .D(
        \fadd_0_0_0_0_4/fracrclose1 [3]), .CLK(clk), .QN(n11901) );
  DFFX1 \fadd_0_0_0_0_4/norm/n351_q_reg[4]  ( .D(
        \fadd_0_0_0_0_4/fracrclose1 [4]), .CLK(clk), .QN(n11900) );
  DFFX1 \fadd_0_0_0_0_4/norm/n351_q_reg[5]  ( .D(
        \fadd_0_0_0_0_4/fracrclose1 [5]), .CLK(clk), .Q(n13544), .QN(n11899)
         );
  DFFX1 \fadd_0_0_0_0_4/norm/n352_q_reg[4]  ( .D(
        \fadd_0_0_0_0_4/norm/level1 [4]), .CLK(clk), .Q(
        \fadd_0_0_0_0_4/norm/level1_d1[4] ) );
  DFFX1 \fadd_0_0_0_0_4/norm/n353_q_reg  ( .D(\fadd_0_0_0_0_4/sub_784/B[0] ), 
        .CLK(clk), .QN(n12857) );
  DFFX1 \fadd_0_0_0_0_4/norm/n352_q_reg[3]  ( .D(
        \fadd_0_0_0_0_4/norm/level1 [3]), .CLK(clk), .Q(n13693) );
  DFFX1 \fadd_0_0_0_0_4/norm/n352_q_reg[2]  ( .D(
        \fadd_0_0_0_0_4/norm/level1 [2]), .CLK(clk), .Q(n13551) );
  DFFX1 \fadd_0_0_0_0_4/norm/n352_q_reg[1]  ( .D(
        \fadd_0_0_0_0_4/norm/level1 [1]), .CLK(clk), .Q(n13483) );
  DFFX1 \fadd_0_0_0_0_4/norm/n352_q_reg[0]  ( .D(
        \fadd_0_0_0_0_4/norm/level1 [0]), .CLK(clk), .Q(n13672) );
  DFFX1 \fadd_0_0_0_0_5/norm/n351_q_reg[0]  ( .D(
        \fadd_0_0_0_0_5/fracrclose1 [0]), .CLK(clk), .QN(n11545) );
  DFFX1 \fadd_0_0_0_0_5/norm/n351_q_reg[1]  ( .D(
        \fadd_0_0_0_0_5/fracrclose1 [1]), .CLK(clk), .QN(n11546) );
  DFFX1 \fadd_0_0_0_0_5/norm/n351_q_reg[2]  ( .D(
        \fadd_0_0_0_0_5/fracrclose1 [2]), .CLK(clk), .Q(n14053), .QN(n11906)
         );
  DFFX1 \fadd_0_0_0_0_5/norm/n351_q_reg[3]  ( .D(
        \fadd_0_0_0_0_5/fracrclose1 [3]), .CLK(clk), .QN(n11905) );
  DFFX1 \fadd_0_0_0_0_5/norm/n351_q_reg[4]  ( .D(
        \fadd_0_0_0_0_5/fracrclose1 [4]), .CLK(clk), .QN(n11904) );
  DFFX1 \fadd_0_0_0_0_5/norm/n351_q_reg[5]  ( .D(
        \fadd_0_0_0_0_5/fracrclose1 [5]), .CLK(clk), .Q(n13543), .QN(n11903)
         );
  DFFX1 \fadd_0_0_0_0_5/norm/n352_q_reg[4]  ( .D(
        \fadd_0_0_0_0_5/norm/level1 [4]), .CLK(clk), .Q(
        \fadd_0_0_0_0_5/norm/level1_d1[4] ) );
  DFFX1 \fadd_0_0_0_0_5/norm/n353_q_reg  ( .D(\fadd_0_0_0_0_5/sub_784/B[0] ), 
        .CLK(clk), .QN(n12859) );
  DFFX1 \fadd_0_0_0_0_5/norm/n352_q_reg[3]  ( .D(
        \fadd_0_0_0_0_5/norm/level1 [3]), .CLK(clk), .Q(n13703) );
  DFFX1 \fadd_0_0_0_0_5/norm/n352_q_reg[2]  ( .D(
        \fadd_0_0_0_0_5/norm/level1 [2]), .CLK(clk), .Q(n13567) );
  DFFX1 \fadd_0_0_0_0_5/norm/n352_q_reg[1]  ( .D(
        \fadd_0_0_0_0_5/norm/level1 [1]), .CLK(clk), .Q(n13490) );
  DFFX1 \fadd_0_0_0_0_5/norm/n352_q_reg[0]  ( .D(
        \fadd_0_0_0_0_5/norm/level1 [0]), .CLK(clk), .Q(n13682) );
  DFFX1 \fadd_0_0_0_0_6/norm/n351_q_reg[0]  ( .D(
        \fadd_0_0_0_0_6/fracrclose1 [0]), .CLK(clk), .QN(n11558) );
  DFFX1 \fadd_0_0_0_0_6/norm/n351_q_reg[1]  ( .D(
        \fadd_0_0_0_0_6/fracrclose1 [1]), .CLK(clk), .QN(n11559) );
  DFFX1 \fadd_0_0_0_0_6/norm/n351_q_reg[2]  ( .D(
        \fadd_0_0_0_0_6/fracrclose1 [2]), .CLK(clk), .Q(n14054), .QN(n11910)
         );
  DFFX1 \fadd_0_0_0_0_6/norm/n351_q_reg[3]  ( .D(
        \fadd_0_0_0_0_6/fracrclose1 [3]), .CLK(clk), .QN(n11909) );
  DFFX1 \fadd_0_0_0_0_6/norm/n351_q_reg[4]  ( .D(
        \fadd_0_0_0_0_6/fracrclose1 [4]), .CLK(clk), .QN(n11908) );
  DFFX1 \fadd_0_0_0_0_6/norm/n351_q_reg[5]  ( .D(
        \fadd_0_0_0_0_6/fracrclose1 [5]), .CLK(clk), .Q(n13542), .QN(n11907)
         );
  DFFX1 \fadd_0_0_0_0_6/norm/n352_q_reg[4]  ( .D(
        \fadd_0_0_0_0_6/norm/level1 [4]), .CLK(clk), .Q(
        \fadd_0_0_0_0_6/norm/level1_d1[4] ) );
  DFFX1 \fadd_0_0_0_0_6/norm/n353_q_reg  ( .D(\fadd_0_0_0_0_6/sub_784/B[0] ), 
        .CLK(clk), .QN(n12861) );
  DFFX1 \fadd_0_0_0_0_6/norm/n352_q_reg[3]  ( .D(
        \fadd_0_0_0_0_6/norm/level1 [3]), .CLK(clk), .Q(n13699) );
  DFFX1 \fadd_0_0_0_0_6/norm/n352_q_reg[2]  ( .D(
        \fadd_0_0_0_0_6/norm/level1 [2]), .CLK(clk), .Q(n13563) );
  DFFX1 \fadd_0_0_0_0_6/norm/n352_q_reg[1]  ( .D(
        \fadd_0_0_0_0_6/norm/level1 [1]), .CLK(clk), .Q(n13486) );
  DFFX1 \fadd_0_0_0_0_6/norm/n352_q_reg[0]  ( .D(
        \fadd_0_0_0_0_6/norm/level1 [0]), .CLK(clk), .Q(n13678) );
  DFFX1 \fadd_0_0_0_0_7/norm/n351_q_reg[0]  ( .D(
        \fadd_0_0_0_0_7/fracrclose1 [0]), .CLK(clk), .QN(n11571) );
  DFFX1 \fadd_0_0_0_0_7/norm/n351_q_reg[1]  ( .D(
        \fadd_0_0_0_0_7/fracrclose1 [1]), .CLK(clk), .QN(n11572) );
  DFFX1 \fadd_0_0_0_0_7/norm/n351_q_reg[2]  ( .D(
        \fadd_0_0_0_0_7/fracrclose1 [2]), .CLK(clk), .Q(n14055), .QN(n11914)
         );
  DFFX1 \fadd_0_0_0_0_7/norm/n351_q_reg[3]  ( .D(
        \fadd_0_0_0_0_7/fracrclose1 [3]), .CLK(clk), .QN(n11913) );
  DFFX1 \fadd_0_0_0_0_7/norm/n351_q_reg[4]  ( .D(
        \fadd_0_0_0_0_7/fracrclose1 [4]), .CLK(clk), .QN(n11912) );
  DFFX1 \fadd_0_0_0_0_7/norm/n351_q_reg[5]  ( .D(
        \fadd_0_0_0_0_7/fracrclose1 [5]), .CLK(clk), .Q(n13541), .QN(n11911)
         );
  DFFX1 \fadd_0_0_0_0_7/norm/n352_q_reg[4]  ( .D(
        \fadd_0_0_0_0_7/norm/level1 [4]), .CLK(clk), .Q(
        \fadd_0_0_0_0_7/norm/level1_d1[4] ) );
  DFFX1 \fadd_0_0_0_0_7/norm/n353_q_reg  ( .D(\fadd_0_0_0_0_7/sub_784/B[0] ), 
        .CLK(clk), .QN(n12863) );
  DFFX1 \fadd_0_0_0_0_7/norm/n352_q_reg[3]  ( .D(
        \fadd_0_0_0_0_7/norm/level1 [3]), .CLK(clk), .Q(n13704) );
  DFFX1 \fadd_0_0_0_0_7/norm/n352_q_reg[2]  ( .D(
        \fadd_0_0_0_0_7/norm/level1 [2]), .CLK(clk), .Q(n13568) );
  DFFX1 \fadd_0_0_0_0_7/norm/n352_q_reg[1]  ( .D(
        \fadd_0_0_0_0_7/norm/level1 [1]), .CLK(clk), .Q(n13491) );
  DFFX1 \fadd_0_0_0_0_7/norm/n352_q_reg[0]  ( .D(
        \fadd_0_0_0_0_7/norm/level1 [0]), .CLK(clk), .Q(n13683) );
  DFFX1 \fadd_0_0_0_0_8/norm/n351_q_reg[0]  ( .D(
        \fadd_0_0_0_0_8/fracrclose1 [0]), .CLK(clk), .QN(n11584) );
  DFFX1 \fadd_0_0_0_0_8/norm/n351_q_reg[1]  ( .D(
        \fadd_0_0_0_0_8/fracrclose1 [1]), .CLK(clk), .QN(n11585) );
  DFFX1 \fadd_0_0_0_0_8/norm/n351_q_reg[2]  ( .D(
        \fadd_0_0_0_0_8/fracrclose1 [2]), .CLK(clk), .Q(n14056), .QN(n11918)
         );
  DFFX1 \fadd_0_0_0_0_8/norm/n351_q_reg[3]  ( .D(
        \fadd_0_0_0_0_8/fracrclose1 [3]), .CLK(clk), .QN(n11917) );
  DFFX1 \fadd_0_0_0_0_8/norm/n351_q_reg[4]  ( .D(
        \fadd_0_0_0_0_8/fracrclose1 [4]), .CLK(clk), .QN(n11916) );
  DFFX1 \fadd_0_0_0_0_8/norm/n351_q_reg[5]  ( .D(
        \fadd_0_0_0_0_8/fracrclose1 [5]), .CLK(clk), .Q(n13540), .QN(n11915)
         );
  DFFX1 \fadd_0_0_0_0_8/norm/n352_q_reg[4]  ( .D(
        \fadd_0_0_0_0_8/norm/level1 [4]), .CLK(clk), .Q(
        \fadd_0_0_0_0_8/norm/level1_d1[4] ) );
  DFFX1 \fadd_0_0_0_0_8/norm/n353_q_reg  ( .D(\fadd_0_0_0_0_8/sub_784/B[0] ), 
        .CLK(clk), .QN(n12865) );
  DFFX1 \fadd_0_0_0_0_8/norm/n352_q_reg[3]  ( .D(
        \fadd_0_0_0_0_8/norm/level1 [3]), .CLK(clk), .Q(n13692) );
  DFFX1 \fadd_0_0_0_0_8/norm/n352_q_reg[2]  ( .D(
        \fadd_0_0_0_0_8/norm/level1 [2]), .CLK(clk), .Q(n13550) );
  DFFX1 \fadd_0_0_0_0_8/norm/n352_q_reg[1]  ( .D(
        \fadd_0_0_0_0_8/norm/level1 [1]), .CLK(clk), .Q(n13482) );
  DFFX1 \fadd_0_0_0_0_8/norm/n352_q_reg[0]  ( .D(
        \fadd_0_0_0_0_8/norm/level1 [0]), .CLK(clk), .Q(n13671) );
  DFFX1 \fadd_0_0_0_0_9/norm/n351_q_reg[0]  ( .D(
        \fadd_0_0_0_0_9/fracrclose1 [0]), .CLK(clk), .QN(n11597) );
  DFFX1 \fadd_0_0_0_0_9/norm/n351_q_reg[1]  ( .D(
        \fadd_0_0_0_0_9/fracrclose1 [1]), .CLK(clk), .QN(n11598) );
  DFFX1 \fadd_0_0_0_0_9/norm/n351_q_reg[2]  ( .D(
        \fadd_0_0_0_0_9/fracrclose1 [2]), .CLK(clk), .Q(n14057), .QN(n11922)
         );
  DFFX1 \fadd_0_0_0_0_9/norm/n351_q_reg[3]  ( .D(
        \fadd_0_0_0_0_9/fracrclose1 [3]), .CLK(clk), .QN(n11921) );
  DFFX1 \fadd_0_0_0_0_9/norm/n351_q_reg[4]  ( .D(
        \fadd_0_0_0_0_9/fracrclose1 [4]), .CLK(clk), .QN(n11920) );
  DFFX1 \fadd_0_0_0_0_9/norm/n351_q_reg[5]  ( .D(
        \fadd_0_0_0_0_9/fracrclose1 [5]), .CLK(clk), .Q(n13539), .QN(n11919)
         );
  DFFX1 \fadd_0_0_0_0_9/norm/n352_q_reg[4]  ( .D(
        \fadd_0_0_0_0_9/norm/level1 [4]), .CLK(clk), .Q(
        \fadd_0_0_0_0_9/norm/level1_d1[4] ) );
  DFFX1 \fadd_0_0_0_0_9/norm/n353_q_reg  ( .D(\fadd_0_0_0_0_9/sub_784/B[0] ), 
        .CLK(clk), .QN(n12867) );
  DFFX1 \fadd_0_0_0_0_9/norm/n352_q_reg[3]  ( .D(
        \fadd_0_0_0_0_9/norm/level1 [3]), .CLK(clk), .Q(n13705) );
  DFFX1 \fadd_0_0_0_0_9/norm/n352_q_reg[2]  ( .D(
        \fadd_0_0_0_0_9/norm/level1 [2]), .CLK(clk), .Q(n13569) );
  DFFX1 \fadd_0_0_0_0_9/norm/n352_q_reg[1]  ( .D(
        \fadd_0_0_0_0_9/norm/level1 [1]), .CLK(clk), .Q(n13492) );
  DFFX1 \fadd_0_0_0_0_9/norm/n352_q_reg[0]  ( .D(
        \fadd_0_0_0_0_9/norm/level1 [0]), .CLK(clk), .Q(n13684) );
  DFFX1 \fmul_0_0_0_0_0/n114_q_reg[0]  ( .D(\fmul_0_0_0_0_0/exc [0]), .CLK(clk), .Q(n11954) );
  DFFX1 \fmul_0_0_0_0_0/n114_q_reg[1]  ( .D(\fmul_0_0_0_0_0/exc [1]), .CLK(clk), .Q(n13754), .QN(n11953) );
  DFFX1 \fmul_0_0_0_0_0/n113_q_reg  ( .D(\fmul_0_0_0_0_0/sign ), .CLK(clk), 
        .Q(\U565/DATA2_9 ) );
  DFFX1 \fmul_0_0_0_0_1/n114_q_reg[0]  ( .D(\fmul_0_0_0_0_1/exc [0]), .CLK(clk), .Q(n13766) );
  DFFX1 \fmul_0_0_0_0_1/n114_q_reg[1]  ( .D(\fmul_0_0_0_0_1/exc [1]), .CLK(clk), .Q(n11939) );
  DFFX1 \fmul_0_0_0_0_1/n113_q_reg  ( .D(\fmul_0_0_0_0_1/sign ), .CLK(clk), 
        .Q(\U503/DATA2_9 ) );
  DFFX1 \fadd_0_0_0_0_1_y_reg[9]  ( .D(n13126), .CLK(clk), .Q(n13717), .QN(
        n11665) );
  DFFX1 \fmul_0_0_0_0_2/n114_q_reg[0]  ( .D(\fmul_0_0_0_0_2/exc [0]), .CLK(clk), .Q(n13751) );
  DFFX1 \fmul_0_0_0_0_2/n114_q_reg[1]  ( .D(\fmul_0_0_0_0_2/exc [1]), .CLK(clk), .Q(n11943), .QN(n13781) );
  DFFX1 \fmul_0_0_0_0_2/n113_q_reg  ( .D(\fmul_0_0_0_0_2/sign ), .CLK(clk), 
        .Q(\U450/DATA2_9 ) );
  DFFX1 \fmul_0_0_0_0_3/n114_q_reg[0]  ( .D(\fmul_0_0_0_0_3/exc [0]), .CLK(clk), .Q(n13767) );
  DFFX1 \fmul_0_0_0_0_3/n114_q_reg[1]  ( .D(\fmul_0_0_0_0_3/exc [1]), .CLK(clk), .Q(n11941) );
  DFFX1 \fmul_0_0_0_0_3/n113_q_reg  ( .D(\fmul_0_0_0_0_3/sign ), .CLK(clk), 
        .Q(\U394/DATA2_9 ) );
  DFFX1 \fadd_0_0_0_0_3_y_reg[9]  ( .D(n13102), .CLK(clk), .Q(n13718), .QN(
        n11686) );
  DFFX1 \fmul_0_0_0_0_4/n114_q_reg[0]  ( .D(\fmul_0_0_0_0_4/exc [0]), .CLK(clk), .Q(n13747) );
  DFFX1 \fmul_0_0_0_0_4/n114_q_reg[1]  ( .D(\fmul_0_0_0_0_4/exc [1]), .CLK(clk), .Q(n11951), .QN(n13750) );
  DFFX1 \fmul_0_0_0_0_4/n113_q_reg  ( .D(\fmul_0_0_0_0_4/sign ), .CLK(clk), 
        .Q(\U341/DATA2_9 ) );
  DFFX1 \fmul_0_0_0_0_5/n114_q_reg[0]  ( .D(\fmul_0_0_0_0_5/exc [0]), .CLK(clk), .Q(n13768) );
  DFFX1 \fmul_0_0_0_0_5/n114_q_reg[1]  ( .D(\fmul_0_0_0_0_5/exc [1]), .CLK(clk), .Q(n11945) );
  DFFX1 \fmul_0_0_0_0_5/n113_q_reg  ( .D(\fmul_0_0_0_0_5/sign ), .CLK(clk), 
        .Q(\U282/DATA2_9 ) );
  DFFX1 \fadd_0_0_0_0_5_y_reg[9]  ( .D(n13054), .CLK(clk), .Q(n13719), .QN(
        n11728) );
  DFFX1 \fmul_0_0_0_0_6/n114_q_reg[0]  ( .D(\fmul_0_0_0_0_6/exc [0]), .CLK(clk), .Q(n13752) );
  DFFX1 \fmul_0_0_0_0_6/n114_q_reg[1]  ( .D(\fmul_0_0_0_0_6/exc [1]), .CLK(clk), .Q(n11949), .QN(n13780) );
  DFFX1 \fmul_0_0_0_0_6/n113_q_reg  ( .D(\fmul_0_0_0_0_6/sign ), .CLK(clk), 
        .Q(\U229/DATA2_9 ) );
  DFFX1 \fmul_0_0_0_0_7/n114_q_reg[0]  ( .D(\fmul_0_0_0_0_7/exc [0]), .CLK(clk), .Q(n13769) );
  DFFX1 \fmul_0_0_0_0_7/n114_q_reg[1]  ( .D(\fmul_0_0_0_0_7/exc [1]), .CLK(clk), .Q(n11947) );
  DFFX1 \fmul_0_0_0_0_7/n113_q_reg  ( .D(\fmul_0_0_0_0_7/sign ), .CLK(clk), 
        .Q(\U173/DATA2_9 ) );
  DFFX1 \fadd_0_0_0_0_7_y_reg[9]  ( .D(n13030), .CLK(clk), .Q(n13720), .QN(
        n11749) );
  DFFX1 \fmul_0_0_0_0_8/n114_q_reg[0]  ( .D(\fmul_0_0_0_0_8/exc [0]), .CLK(clk), .Q(n13753), .QN(n11960) );
  DFFX1 \fmul_0_0_0_0_8/n114_q_reg[1]  ( .D(\fmul_0_0_0_0_8/exc [1]), .CLK(clk), .Q(n11961) );
  DFFX1 \fmul_0_0_0_0_8/n113_q_reg  ( .D(\fmul_0_0_0_0_8/sign ), .CLK(clk), 
        .QN(n11866) );
  DFFX1 \fmul_0_0_0_0_9/n114_q_reg[0]  ( .D(\fmul_0_0_0_0_9/exc [0]), .CLK(clk), .Q(n13770) );
  DFFX1 \fmul_0_0_0_0_9/n114_q_reg[1]  ( .D(\fmul_0_0_0_0_9/exc [1]), .CLK(clk), .Q(n11956) );
  DFFX1 \fmul_0_0_0_0_9/n113_q_reg  ( .D(\fmul_0_0_0_0_9/sign ), .CLK(clk), 
        .Q(\U58/DATA2_9 ) );
  DFFX1 \fadd_0_0_0_0_9_y_reg[9]  ( .D(n12934), .CLK(clk), .Q(n13721), .QN(
        n11833) );
  DFFX1 \fmul_0_0_0_0_10/n114_q_reg[0]  ( .D(\fmul_0_0_0_0_10/U9/Z_0 ), .CLK(
        clk), .Q(n13771) );
  DFFX1 \fmul_0_0_0_0_10/n114_q_reg[1]  ( .D(\fmul_0_0_0_0_10/U9/Z_1 ), .CLK(
        clk), .Q(n11958) );
  DFFX1 \fmul_0_0_0_0_10/n113_q_reg  ( .D(\fmul_0_0_0_0_10/n137 ), .CLK(clk), 
        .Q(\U5/DATA2_9 ) );
  DFFX1 \fadd_0_0_0_0_10_y_reg[9]  ( .D(n12910), .CLK(clk), .Q(n13726), .QN(
        n11849) );
  DFFX1 \fmul_0_0_0_0_0/roundingadder/n155_q_reg[0]  ( .D(
        \fmul_0_0_0_0_0/sigprodext [6]), .CLK(clk), .Q(
        \fmul_0_0_0_0_0/roundingadder/x_1_d1 [0]) );
  DFFX1 \fmul_0_0_0_0_0/roundingadder/n155_q_reg[1]  ( .D(
        \fmul_0_0_0_0_0/sigprodext [7]), .CLK(clk), .Q(
        \fmul_0_0_0_0_0/roundingadder/x_1_d1 [1]) );
  DFFX1 \fmul_0_0_0_0_0/roundingadder/n155_q_reg[2]  ( .D(
        \fmul_0_0_0_0_0/sigprodext [8]), .CLK(clk), .Q(
        \fmul_0_0_0_0_0/roundingadder/x_1_d1 [2]) );
  DFFX1 \fmul_0_0_0_0_0/roundingadder/n155_q_reg[3]  ( .D(
        \fmul_0_0_0_0_0/sigprodext [9]), .CLK(clk), .Q(
        \fmul_0_0_0_0_0/roundingadder/x_1_d1 [3]) );
  DFFX1 \fmul_0_0_0_0_0/roundingadder/n155_q_reg[4]  ( .D(
        \fmul_0_0_0_0_0/exppostnorm [0]), .CLK(clk), .Q(
        \fmul_0_0_0_0_0/roundingadder/x_1_d1 [4]) );
  DFFX1 \fmul_0_0_0_0_0/roundingadder/n155_q_reg[5]  ( .D(
        \fmul_0_0_0_0_0/exppostnorm [1]), .CLK(clk), .Q(
        \fmul_0_0_0_0_0/roundingadder/x_1_d1 [5]) );
  DFFX1 \fmul_0_0_0_0_0/roundingadder/n155_q_reg[6]  ( .D(
        \fmul_0_0_0_0_0/exppostnorm [2]), .CLK(clk), .Q(
        \fmul_0_0_0_0_0/roundingadder/x_1_d1 [6]) );
  DFFX1 \fmul_0_0_0_0_0/roundingadder/n155_q_reg[7]  ( .D(
        \fmul_0_0_0_0_0/exppostnorm [3]), .CLK(clk), .Q(
        \fmul_0_0_0_0_0/roundingadder/x_1_d1 [7]) );
  DFFX1 \fmul_0_0_0_0_0/roundingadder/n155_q_reg[8]  ( .D(
        \fmul_0_0_0_0_0/exppostnorm [4]), .CLK(clk), .Q(
        \fmul_0_0_0_0_0/roundingadder/x_1_d1 [8]) );
  DFFX1 \fmul_0_0_0_0_0/roundingadder/n155_q_reg[9]  ( .D(
        \fmul_0_0_0_0_0/exppostnorm [5]), .CLK(clk), .Q(
        \fmul_0_0_0_0_0/roundingadder/x_1_d1 [9]) );
  DFFX1 \fmul_0_0_0_0_0/roundingadder/n155_q_reg[10]  ( .D(n14127), .CLK(clk), 
        .Q(\fmul_0_0_0_0_0/roundingadder/x_1_d1 [10]) );
  DFFX1 \fmul_0_0_0_0_0/roundingadder/n154_q_reg  ( .D(\fmul_0_0_0_0_0/round ), 
        .CLK(clk), .Q(\fmul_0_0_0_0_0/roundingadder/n151_o[0] ) );
  DFFX1 \fmul_0_0_0_0_1/roundingadder/n155_q_reg[0]  ( .D(
        \fmul_0_0_0_0_1/sigprodext [6]), .CLK(clk), .Q(
        \fmul_0_0_0_0_1/roundingadder/x_1_d1 [0]) );
  DFFX1 \fmul_0_0_0_0_1/roundingadder/n155_q_reg[1]  ( .D(
        \fmul_0_0_0_0_1/sigprodext [7]), .CLK(clk), .Q(
        \fmul_0_0_0_0_1/roundingadder/x_1_d1 [1]) );
  DFFX1 \fmul_0_0_0_0_1/roundingadder/n155_q_reg[2]  ( .D(
        \fmul_0_0_0_0_1/sigprodext [8]), .CLK(clk), .Q(
        \fmul_0_0_0_0_1/roundingadder/x_1_d1 [2]) );
  DFFX1 \fmul_0_0_0_0_1/roundingadder/n155_q_reg[3]  ( .D(
        \fmul_0_0_0_0_1/sigprodext [9]), .CLK(clk), .Q(
        \fmul_0_0_0_0_1/roundingadder/x_1_d1 [3]) );
  DFFX1 \fmul_0_0_0_0_1/roundingadder/n155_q_reg[4]  ( .D(
        \fmul_0_0_0_0_1/exppostnorm [0]), .CLK(clk), .Q(
        \fmul_0_0_0_0_1/roundingadder/x_1_d1 [4]) );
  DFFX1 \fmul_0_0_0_0_1/roundingadder/n155_q_reg[5]  ( .D(
        \fmul_0_0_0_0_1/exppostnorm [1]), .CLK(clk), .Q(
        \fmul_0_0_0_0_1/roundingadder/x_1_d1 [5]) );
  DFFX1 \fmul_0_0_0_0_1/roundingadder/n155_q_reg[6]  ( .D(
        \fmul_0_0_0_0_1/exppostnorm [2]), .CLK(clk), .Q(
        \fmul_0_0_0_0_1/roundingadder/x_1_d1 [6]) );
  DFFX1 \fmul_0_0_0_0_1/roundingadder/n155_q_reg[7]  ( .D(
        \fmul_0_0_0_0_1/exppostnorm [3]), .CLK(clk), .Q(
        \fmul_0_0_0_0_1/roundingadder/x_1_d1 [7]) );
  DFFX1 \fmul_0_0_0_0_1/roundingadder/n155_q_reg[8]  ( .D(
        \fmul_0_0_0_0_1/exppostnorm [4]), .CLK(clk), .Q(
        \fmul_0_0_0_0_1/roundingadder/x_1_d1 [8]) );
  DFFX1 \fmul_0_0_0_0_1/roundingadder/n155_q_reg[9]  ( .D(
        \fmul_0_0_0_0_1/exppostnorm [5]), .CLK(clk), .Q(
        \fmul_0_0_0_0_1/roundingadder/x_1_d1 [9]) );
  DFFX1 \fmul_0_0_0_0_1/roundingadder/n155_q_reg[10]  ( .D(n14136), .CLK(clk), 
        .Q(\fmul_0_0_0_0_1/roundingadder/x_1_d1 [10]) );
  DFFX1 \fmul_0_0_0_0_1/roundingadder/n154_q_reg  ( .D(\fmul_0_0_0_0_1/round ), 
        .CLK(clk), .Q(\fmul_0_0_0_0_1/roundingadder/n151_o[0] ) );
  DFFX1 \fadd_0_0_0_0_1_y_reg[0]  ( .D(n13135), .CLK(clk), .Q(n13637), .QN(
        n11656) );
  DFFX1 \fadd_0_0_0_0_1_y_reg[1]  ( .D(n13134), .CLK(clk), .Q(n13665), .QN(
        n11657) );
  DFFX1 \fadd_0_0_0_0_1_y_reg[2]  ( .D(n13133), .CLK(clk), .Q(n13686), .QN(
        n11658) );
  DFFX1 \fadd_0_0_0_0_1_y_reg[3]  ( .D(n13132), .CLK(clk), .Q(n13708), .QN(
        n11659) );
  DFFX1 \fadd_0_0_0_0_1_y_reg[4]  ( .D(n13131), .CLK(clk), .Q(n5910), .QN(
        n14546) );
  DFFX1 \fadd_0_0_0_0_1_y_reg[5]  ( .D(n13130), .CLK(clk), .Q(n5911), .QN(
        n14545) );
  DFFX1 \fadd_0_0_0_0_1_y_reg[6]  ( .D(n13129), .CLK(clk), .Q(n5912), .QN(
        n14544) );
  DFFX1 \fadd_0_0_0_0_1_y_reg[7]  ( .D(n13128), .CLK(clk), .Q(n5913), .QN(
        n14543) );
  DFFX1 \fadd_0_0_0_0_1_y_reg[8]  ( .D(n13127), .CLK(clk), .Q(n5914), .QN(
        n14542) );
  DFFX1 \fadd_0_0_0_0_1_y_reg[11]  ( .D(n13124), .CLK(clk), .Q(n13622), .QN(
        n12706) );
  DFFX1 \fadd_0_0_0_0_1_y_reg[10]  ( .D(n13125), .CLK(clk), .Q(n13889), .QN(
        n11666) );
  DFFX1 \fadd_0_0_0_0_1/n293_q_reg[0]  ( .D(\fadd_0_0_0_0_1/newy_10 ), .CLK(
        clk), .Q(\fadd_0_0_0_0_1/syncexnxy_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_1/n294_q_reg[0]  ( .D(\fadd_0_0_0_0_1/syncexnxy_d1 [0]), 
        .CLK(clk), .Q(n12361) );
  DFFX1 \p_val_59_reg[9]  ( .D(n12688), .CLK(clk), .Q(n13968) );
  DFFX1 \p_val_288_reg[9]  ( .D(n12687), .CLK(clk), .Q(n13811) );
  DFFX1 \fadd_0_0_0_0_1_x_reg[9]  ( .D(n13114), .CLK(clk), .Q(n13579), .QN(
        n11676) );
  DFFX1 \fadd_0_0_0_0_1/n288_q_reg  ( .D(\fadd_0_0_0_0_1/newy_9 ), .CLK(clk), 
        .Q(\fadd_0_0_0_0_1/syncsigny_d1 ) );
  DFFX1 \fadd_0_0_0_0_1/n289_q_reg  ( .D(\fadd_0_0_0_0_1/syncsigny_d1 ), .CLK(
        clk), .QN(n12358) );
  DFFX1 \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[7]  ( .D(
        n12702), .CLK(clk), .Q(
        \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [7]) );
  DFFX1 \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[7]  ( .D(
        \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [7]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [7]) );
  DFFX1 \fadd_0_0_0_0_1/n284_q_reg  ( .D(n12702), .CLK(clk), .Q(
        \fadd_0_0_0_0_1/synceffsub_d1 ) );
  DFFX1 \fadd_0_0_0_0_1/n285_q_reg  ( .D(\fadd_0_0_0_0_1/synceffsub_d1 ), 
        .CLK(clk), .QN(n12351) );
  DFFX1 \fadd_0_0_0_0_1/n276_q_reg  ( .D(n12702), .CLK(clk), .Q(
        \fadd_0_0_0_0_1/effsub_d1 ) );
  DFFX1 \fadd_0_0_0_0_1/n277_q_reg  ( .D(\fadd_0_0_0_0_1/effsub_d1 ), .CLK(clk), .QN(n11483) );
  DFFX1 \p_val_59_reg[11]  ( .D(n12686), .CLK(clk), .Q(n13969) );
  DFFX1 \p_val_288_reg[11]  ( .D(n12685), .CLK(clk), .Q(n13812) );
  DFFX1 \fadd_0_0_0_0_1_x_reg[11]  ( .D(n13112), .CLK(clk), .Q(n13509), .QN(
        n12704) );
  DFFX1 \fadd_0_0_0_0_1/n293_q_reg[3]  ( .D(\fadd_0_0_0_0_1/newx [11]), .CLK(
        clk), .Q(\fadd_0_0_0_0_1/syncexnxy_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_1/n294_q_reg[3]  ( .D(\fadd_0_0_0_0_1/syncexnxy_d1 [3]), 
        .CLK(clk), .Q(n13774), .QN(n12359) );
  DFFX1 \p_val_59_reg[10]  ( .D(n12684), .CLK(clk), .Q(n13970) );
  DFFX1 \p_val_288_reg[10]  ( .D(n12683), .CLK(clk), .Q(n13813) );
  DFFX1 \fadd_0_0_0_0_1_x_reg[10]  ( .D(n13113), .CLK(clk), .Q(n13502), .QN(
        n12705) );
  DFFX1 \fadd_0_0_0_0_1/n286_q_reg[9]  ( .D(n14679), .CLK(clk), .Q(
        \fadd_0_0_0_0_1/syncx_d1 [9]) );
  DFFX1 \fadd_0_0_0_0_1/n287_q_reg[9]  ( .D(\fadd_0_0_0_0_1/syncx_d1 [9]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_1/syncx_d2 [9]) );
  DFFX1 \fadd_0_0_0_0_1/n286_q_reg[0]  ( .D(
        \add_0_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .CLK(clk), .Q(\fadd_0_0_0_0_1/syncx_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_1/n287_q_reg[0]  ( .D(\fadd_0_0_0_0_1/syncx_d1 [0]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_1/syncx_d2 [0]) );
  DFFX1 \p_val_59_reg[0]  ( .D(n12682), .CLK(clk), .Q(n13971) );
  DFFX1 \p_val_288_reg[0]  ( .D(n12681), .CLK(clk), .Q(n14082), .QN(n12348) );
  DFFX1 \fadd_0_0_0_0_1_x_reg[0]  ( .D(n13123), .CLK(clk), .Q(n13517), .QN(
        n11667) );
  DFFX1 \fadd_0_0_0_0_1/rightshiftercomponent/n415_q_reg[2]  ( .D(n14683), 
        .CLK(clk), .QN(n11489) );
  DFFX1 \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/n432_q_reg[2]  ( .D(
        \add_0_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .CLK(clk), .Q(\fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/n433_q_reg[2]  ( .D(
        \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [2]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/x_d2 [2]) );
  DFFX1 \fadd_0_0_0_0_1/n293_q_reg[2]  ( .D(\fadd_0_0_0_0_1/newx [10]), .CLK(
        clk), .Q(\fadd_0_0_0_0_1/syncexnxy_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_1/n294_q_reg[2]  ( .D(\fadd_0_0_0_0_1/syncexnxy_d1 [2]), 
        .CLK(clk), .Q(n13730), .QN(n12357) );
  DFFX1 \fadd_0_0_0_0_1/n286_q_reg[1]  ( .D(
        \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ), .CLK(clk), .Q(\fadd_0_0_0_0_1/syncx_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_1/n287_q_reg[1]  ( .D(\fadd_0_0_0_0_1/syncx_d1 [1]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_1/syncx_d2 [1]) );
  DFFX1 \p_val_59_reg[1]  ( .D(n12680), .CLK(clk), .Q(n13972) );
  DFFX1 \p_val_288_reg[1]  ( .D(n12679), .CLK(clk), .Q(n14083), .QN(n12346) );
  DFFX1 \fadd_0_0_0_0_1_x_reg[1]  ( .D(n13122), .CLK(clk), .Q(n13528), .QN(
        n11668) );
  DFFX1 \fadd_0_0_0_0_1/rightshiftercomponent/n415_q_reg[3]  ( .D(n14682), 
        .CLK(clk), .QN(n11490) );
  DFFX1 \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/n432_q_reg[3]  ( .D(
        \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ), .CLK(clk), .Q(\fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/n433_q_reg[3]  ( .D(
        \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [3]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/x_d2 [3]) );
  DFFX1 \fadd_0_0_0_0_1/n286_q_reg[2]  ( .D(
        \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ), .CLK(clk), .Q(\fadd_0_0_0_0_1/syncx_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_1/n287_q_reg[2]  ( .D(\fadd_0_0_0_0_1/syncx_d1 [2]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_1/syncx_d2 [2]) );
  DFFX1 \p_val_59_reg[2]  ( .D(n12678), .CLK(clk), .Q(n13973) );
  DFFX1 \p_val_288_reg[2]  ( .D(n12677), .CLK(clk), .Q(n14084), .QN(n12344) );
  DFFX1 \fadd_0_0_0_0_1_x_reg[2]  ( .D(n13121), .CLK(clk), .Q(n13553), .QN(
        n11669) );
  DFFX1 \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/n432_q_reg[4]  ( .D(
        \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ), .CLK(clk), .Q(\fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/n433_q_reg[4]  ( .D(
        \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [4]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/x_d2 [4]) );
  DFFX1 \fadd_0_0_0_0_1/n286_q_reg[3]  ( .D(
        \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ), .CLK(clk), .Q(\fadd_0_0_0_0_1/syncx_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_1/n287_q_reg[3]  ( .D(\fadd_0_0_0_0_1/syncx_d1 [3]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_1/syncx_d2 [3]) );
  DFFX1 \p_val_59_reg[3]  ( .D(n12676), .CLK(clk), .Q(n13974) );
  DFFX1 \p_val_288_reg[3]  ( .D(n12675), .CLK(clk), .Q(n14085), .QN(n12342) );
  DFFX1 \fadd_0_0_0_0_1_x_reg[3]  ( .D(n13120), .CLK(clk), .Q(n13570), .QN(
        n11670) );
  DFFX1 \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/n432_q_reg[5]  ( .D(
        \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ), .CLK(clk), .Q(\fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [5]) );
  DFFX1 \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/n433_q_reg[5]  ( .D(
        \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [5]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/x_d2 [5]) );
  DFFX1 \fadd_0_0_0_0_1/n275_q_reg[4]  ( .D(\fadd_0_0_0_0_1/newx [4]), .CLK(
        clk), .Q(\fadd_0_0_0_0_1/newx_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_1/n281_q_reg[0]  ( .D(\fadd_0_0_0_0_1/newx [4]), .CLK(
        clk), .Q(\fadd_0_0_0_0_1/exponentresultfar0_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_1/n282_q_reg[0]  ( .D(
        \fadd_0_0_0_0_1/exponentresultfar0_d1 [0]), .CLK(clk), .Q(
        \fadd_0_0_0_0_1/exponentresultfar0_d2 [0]) );
  DFFX1 \fadd_0_0_0_0_1/n286_q_reg[4]  ( .D(\fadd_0_0_0_0_1/newx [4]), .CLK(
        clk), .Q(\fadd_0_0_0_0_1/syncx_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_1/n287_q_reg[4]  ( .D(\fadd_0_0_0_0_1/syncx_d1 [4]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_1/syncx_d2 [4]) );
  DFFX1 \p_val_59_reg[4]  ( .D(n12674), .CLK(clk), .Q(n13975) );
  DFFX1 \p_val_288_reg[4]  ( .D(n12673), .CLK(clk), .Q(n14086), .QN(n12340) );
  DFFX1 \fadd_0_0_0_0_1_x_reg[4]  ( .D(n13119), .CLK(clk), .Q(n5922), .QN(
        n14551) );
  DFFX1 \fadd_0_0_0_0_1/n275_q_reg[5]  ( .D(\fadd_0_0_0_0_1/newx [5]), .CLK(
        clk), .Q(\fadd_0_0_0_0_1/newx_d1 [5]) );
  DFFX1 \fadd_0_0_0_0_1/n281_q_reg[1]  ( .D(\fadd_0_0_0_0_1/newx [5]), .CLK(
        clk), .Q(\fadd_0_0_0_0_1/exponentresultfar0_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_1/n282_q_reg[1]  ( .D(
        \fadd_0_0_0_0_1/exponentresultfar0_d1 [1]), .CLK(clk), .Q(
        \fadd_0_0_0_0_1/exponentresultfar0_d2 [1]) );
  DFFX1 \fadd_0_0_0_0_1/n286_q_reg[5]  ( .D(\fadd_0_0_0_0_1/newx [5]), .CLK(
        clk), .Q(\fadd_0_0_0_0_1/syncx_d1 [5]) );
  DFFX1 \fadd_0_0_0_0_1/n287_q_reg[5]  ( .D(\fadd_0_0_0_0_1/syncx_d1 [5]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_1/syncx_d2 [5]) );
  DFFX1 \p_val_59_reg[5]  ( .D(n12672), .CLK(clk), .Q(n13976) );
  DFFX1 \p_val_288_reg[5]  ( .D(n12671), .CLK(clk), .Q(n14087), .QN(n12338) );
  DFFX1 \fadd_0_0_0_0_1_x_reg[5]  ( .D(n13118), .CLK(clk), .Q(n5923), .QN(
        n14550) );
  DFFX1 \fadd_0_0_0_0_1/n275_q_reg[6]  ( .D(\fadd_0_0_0_0_1/newx [6]), .CLK(
        clk), .Q(\fadd_0_0_0_0_1/newx_d1 [6]) );
  DFFX1 \fadd_0_0_0_0_1/n281_q_reg[2]  ( .D(\fadd_0_0_0_0_1/newx [6]), .CLK(
        clk), .Q(\fadd_0_0_0_0_1/exponentresultfar0_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_1/n282_q_reg[2]  ( .D(
        \fadd_0_0_0_0_1/exponentresultfar0_d1 [2]), .CLK(clk), .Q(
        \fadd_0_0_0_0_1/exponentresultfar0_d2 [2]) );
  DFFX1 \fadd_0_0_0_0_1/n286_q_reg[6]  ( .D(\fadd_0_0_0_0_1/newx [6]), .CLK(
        clk), .Q(\fadd_0_0_0_0_1/syncx_d1 [6]) );
  DFFX1 \fadd_0_0_0_0_1/n287_q_reg[6]  ( .D(\fadd_0_0_0_0_1/syncx_d1 [6]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_1/syncx_d2 [6]) );
  DFFX1 \p_val_59_reg[6]  ( .D(n12670), .CLK(clk), .Q(n13977) );
  DFFX1 \p_val_288_reg[6]  ( .D(n12669), .CLK(clk), .Q(n14088), .QN(n12336) );
  DFFX1 \fadd_0_0_0_0_1_x_reg[6]  ( .D(n13117), .CLK(clk), .Q(n5924), .QN(
        n14549) );
  DFFX1 \fadd_0_0_0_0_1/n275_q_reg[7]  ( .D(\fadd_0_0_0_0_1/newx [7]), .CLK(
        clk), .Q(\fadd_0_0_0_0_1/newx_d1 [7]) );
  DFFX1 \fadd_0_0_0_0_1/n281_q_reg[3]  ( .D(\fadd_0_0_0_0_1/newx [7]), .CLK(
        clk), .Q(\fadd_0_0_0_0_1/exponentresultfar0_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_1/n282_q_reg[3]  ( .D(
        \fadd_0_0_0_0_1/exponentresultfar0_d1 [3]), .CLK(clk), .Q(
        \fadd_0_0_0_0_1/exponentresultfar0_d2 [3]) );
  DFFX1 \fadd_0_0_0_0_1/n286_q_reg[7]  ( .D(\fadd_0_0_0_0_1/newx [7]), .CLK(
        clk), .Q(\fadd_0_0_0_0_1/syncx_d1 [7]) );
  DFFX1 \fadd_0_0_0_0_1/n287_q_reg[7]  ( .D(\fadd_0_0_0_0_1/syncx_d1 [7]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_1/syncx_d2 [7]) );
  DFFX1 \p_val_59_reg[7]  ( .D(n12668), .CLK(clk), .Q(n13978) );
  DFFX1 \p_val_288_reg[7]  ( .D(n12667), .CLK(clk), .Q(n14089), .QN(n12334) );
  DFFX1 \fadd_0_0_0_0_1_x_reg[7]  ( .D(n13116), .CLK(clk), .Q(n5925), .QN(
        n14548) );
  DFFX1 \fadd_0_0_0_0_1/n275_q_reg[8]  ( .D(\fadd_0_0_0_0_1/newx [8]), .CLK(
        clk), .Q(\fadd_0_0_0_0_1/newx_d1 [8]) );
  DFFX1 \fadd_0_0_0_0_1/n280_q_reg[0]  ( .D(
        \fadd_0_0_0_0_1/exponentresultclose [0]), .CLK(clk), .Q(
        \fadd_0_0_0_0_1/exponentresultclose_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_1/n280_q_reg[1]  ( .D(
        \fadd_0_0_0_0_1/exponentresultclose [1]), .CLK(clk), .Q(
        \fadd_0_0_0_0_1/exponentresultclose_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_1/n280_q_reg[2]  ( .D(
        \fadd_0_0_0_0_1/exponentresultclose [2]), .CLK(clk), .Q(
        \fadd_0_0_0_0_1/exponentresultclose_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_1/n280_q_reg[3]  ( .D(
        \fadd_0_0_0_0_1/exponentresultclose [3]), .CLK(clk), .Q(
        \fadd_0_0_0_0_1/exponentresultclose_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_1/n280_q_reg[4]  ( .D(
        \fadd_0_0_0_0_1/exponentresultclose [4]), .CLK(clk), .Q(
        \fadd_0_0_0_0_1/exponentresultclose_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_1/n280_q_reg[6]  ( .D(n13663), .CLK(clk), .Q(
        \fadd_0_0_0_0_1/exponentresultclose_d1 [6]) );
  DFFX1 \fadd_0_0_0_0_1/n280_q_reg[5]  ( .D(n13663), .CLK(clk), .Q(
        \fadd_0_0_0_0_1/exponentresultclose_d1 [5]) );
  DFFX1 \fadd_0_0_0_0_1/n281_q_reg[4]  ( .D(\fadd_0_0_0_0_1/newx [8]), .CLK(
        clk), .Q(\fadd_0_0_0_0_1/exponentresultfar0_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_1/n282_q_reg[4]  ( .D(
        \fadd_0_0_0_0_1/exponentresultfar0_d1 [4]), .CLK(clk), .Q(
        \fadd_0_0_0_0_1/exponentresultfar0_d2 [4]) );
  DFFX1 \fadd_0_0_0_0_1/n286_q_reg[8]  ( .D(\fadd_0_0_0_0_1/newx [8]), .CLK(
        clk), .Q(\fadd_0_0_0_0_1/syncx_d1 [8]) );
  DFFX1 \fadd_0_0_0_0_1/n287_q_reg[8]  ( .D(\fadd_0_0_0_0_1/syncx_d1 [8]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_1/syncx_d2 [8]) );
  DFFX1 \p_val_59_reg[8]  ( .D(n12666), .CLK(clk), .Q(n13979) );
  DFFX1 \p_val_288_reg[8]  ( .D(n12665), .CLK(clk), .Q(n14090), .QN(n12332) );
  DFFX1 \fadd_0_0_0_0_1_x_reg[8]  ( .D(n13115), .CLK(clk), .Q(n5926), .QN(
        n14547) );
  DFFX1 \fadd_0_0_0_0_1/rightshiftercomponent/n413_q_reg[2]  ( .D(n14673), 
        .CLK(clk), .Q(\fadd_0_0_0_0_1/rightshiftercomponent/ps_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_1/rightshiftercomponent/n416_q_reg[1]  ( .D(
        \fadd_0_0_0_0_1/rightshiftercomponent/level2[1] ), .CLK(clk), .QN(
        n11491) );
  DFFX1 \fadd_0_0_0_0_1/rightshiftercomponent/n416_q_reg[0]  ( .D(n12701), 
        .CLK(clk), .QN(n11492) );
  DFFX1 \fadd_0_0_0_0_1/rightshiftercomponent/n413_q_reg[1]  ( .D(n14676), 
        .CLK(clk), .Q(\fadd_0_0_0_0_1/rightshiftercomponent/ps_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_1/rightshiftercomponent/n417_q_reg  ( .D(
        \fadd_0_0_0_0_1/rightshiftercomponent/n389_o ), .CLK(clk), .Q(n14942)
         );
  DFFX1 \fadd_0_0_0_0_1/rightshiftercomponent/n418_q_reg[0]  ( .D(n12700), 
        .CLK(clk), .Q(\fadd_0_0_0_0_1/rightshiftercomponent/level1_d1[0] ) );
  DFFX1 \fadd_0_0_0_0_1/rightshiftercomponent/n419_q_reg[0]  ( .D(
        \fadd_0_0_0_0_1/rightshiftercomponent/level1_d1[0] ), .CLK(clk), .Q(
        \fadd_0_0_0_0_1/rightshiftercomponent/level1_d2[0] ) );
  DFFX1 \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[5]  ( .D(
        \fadd_0_0_0_0_1/fracyfarxorop [5]), .CLK(clk), .Q(
        \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [5]) );
  DFFX1 \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[5]  ( .D(
        \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [5]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [5]) );
  DFFX1 \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[3]  ( .D(
        \fadd_0_0_0_0_1/fracyfarxorop [3]), .CLK(clk), .Q(
        \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[3]  ( .D(
        \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [3]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [3]) );
  DFFX1 \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[2]  ( .D(
        \fadd_0_0_0_0_1/fracyfarxorop [2]), .CLK(clk), .Q(
        \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[2]  ( .D(
        \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [2]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [2]) );
  DFFX1 \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[1]  ( .D(
        \fadd_0_0_0_0_1/fracyfarxorop [1]), .CLK(clk), .Q(
        \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[1]  ( .D(
        \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [1]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [1]) );
  DFFX1 \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[0]  ( .D(
        \fadd_0_0_0_0_1/fracyfarxorop [0]), .CLK(clk), .Q(
        \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[0]  ( .D(
        \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [0]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [0]) );
  DFFX1 \fadd_0_0_0_0_1/rightshiftercomponent/n413_q_reg[0]  ( .D(n12699), 
        .CLK(clk), .Q(\fadd_0_0_0_0_1/rightshiftercomponent/ps_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_1/rightshiftercomponent/n414_q_reg[0]  ( .D(
        \fadd_0_0_0_0_1/rightshiftercomponent/ps_d1 [0]), .CLK(clk), .Q(
        \fadd_0_0_0_0_1/rightshiftercomponent/ps_d2[0] ) );
  DFFX1 \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[4]  ( .D(
        \fadd_0_0_0_0_1/fracyfarxorop [4]), .CLK(clk), .Q(
        \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[4]  ( .D(
        \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [4]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [4]) );
  DFFX1 \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[6]  ( .D(
        \fadd_0_0_0_0_1/fracyfarxorop [6]), .CLK(clk), .Q(
        \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [6]) );
  DFFX1 \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[6]  ( .D(
        \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [6]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [6]) );
  DFFX1 \fadd_0_0_0_0_1/n293_q_reg[1]  ( .D(\fadd_0_0_0_0_1/newy_11 ), .CLK(
        clk), .Q(\fadd_0_0_0_0_1/syncexnxy_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_1/n294_q_reg[1]  ( .D(\fadd_0_0_0_0_1/syncexnxy_d1 [1]), 
        .CLK(clk), .Q(n13741), .QN(n12360) );
  DFFX1 \fadd_0_0_0_0_1/n278_q_reg  ( .D(n14672), .CLK(clk), .Q(
        \fadd_0_0_0_0_1/selectclosepath_d1 ), .QN(n11494) );
  DFFX1 \fadd_0_0_0_0_1/n283_q_reg  ( .D(\fadd_0_0_0_0_1/zerofromclose ), 
        .CLK(clk), .Q(\fadd_0_0_0_0_1/zerofromclose_d1 ) );
  DFFX1 \fadd_0_0_0_0_1/n290_q_reg  ( .D(\fadd_0_0_0_0_1/ressign ), .CLK(clk), 
        .Q(\fadd_0_0_0_0_1/syncressign_d1 ) );
  DFFX1 \fadd_0_0_0_0_1/n291_q_reg  ( .D(\fadd_0_0_0_0_1/syncressign_d1 ), 
        .CLK(clk), .QN(n12362) );
  DFFX1 \fmul_0_0_0_0_2/roundingadder/n155_q_reg[0]  ( .D(
        \fmul_0_0_0_0_2/sigprodext [6]), .CLK(clk), .Q(
        \fmul_0_0_0_0_2/roundingadder/x_1_d1 [0]) );
  DFFX1 \fmul_0_0_0_0_2/roundingadder/n155_q_reg[1]  ( .D(
        \fmul_0_0_0_0_2/sigprodext [7]), .CLK(clk), .Q(
        \fmul_0_0_0_0_2/roundingadder/x_1_d1 [1]) );
  DFFX1 \fmul_0_0_0_0_2/roundingadder/n155_q_reg[2]  ( .D(
        \fmul_0_0_0_0_2/sigprodext [8]), .CLK(clk), .Q(
        \fmul_0_0_0_0_2/roundingadder/x_1_d1 [2]) );
  DFFX1 \fmul_0_0_0_0_2/roundingadder/n155_q_reg[3]  ( .D(
        \fmul_0_0_0_0_2/sigprodext [9]), .CLK(clk), .Q(
        \fmul_0_0_0_0_2/roundingadder/x_1_d1 [3]) );
  DFFX1 \fmul_0_0_0_0_2/roundingadder/n155_q_reg[4]  ( .D(
        \fmul_0_0_0_0_2/exppostnorm [0]), .CLK(clk), .Q(
        \fmul_0_0_0_0_2/roundingadder/x_1_d1 [4]) );
  DFFX1 \fmul_0_0_0_0_2/roundingadder/n155_q_reg[5]  ( .D(
        \fmul_0_0_0_0_2/exppostnorm [1]), .CLK(clk), .Q(
        \fmul_0_0_0_0_2/roundingadder/x_1_d1 [5]) );
  DFFX1 \fmul_0_0_0_0_2/roundingadder/n155_q_reg[6]  ( .D(
        \fmul_0_0_0_0_2/exppostnorm [2]), .CLK(clk), .Q(
        \fmul_0_0_0_0_2/roundingadder/x_1_d1 [6]) );
  DFFX1 \fmul_0_0_0_0_2/roundingadder/n155_q_reg[7]  ( .D(
        \fmul_0_0_0_0_2/exppostnorm [3]), .CLK(clk), .Q(
        \fmul_0_0_0_0_2/roundingadder/x_1_d1 [7]) );
  DFFX1 \fmul_0_0_0_0_2/roundingadder/n155_q_reg[8]  ( .D(
        \fmul_0_0_0_0_2/exppostnorm [4]), .CLK(clk), .Q(
        \fmul_0_0_0_0_2/roundingadder/x_1_d1 [8]) );
  DFFX1 \fmul_0_0_0_0_2/roundingadder/n155_q_reg[9]  ( .D(
        \fmul_0_0_0_0_2/exppostnorm [5]), .CLK(clk), .Q(
        \fmul_0_0_0_0_2/roundingadder/x_1_d1 [9]) );
  DFFX1 \fmul_0_0_0_0_2/roundingadder/n155_q_reg[10]  ( .D(n14135), .CLK(clk), 
        .Q(\fmul_0_0_0_0_2/roundingadder/x_1_d1 [10]) );
  DFFX1 \fmul_0_0_0_0_2/roundingadder/n154_q_reg  ( .D(\fmul_0_0_0_0_2/round ), 
        .CLK(clk), .Q(\fmul_0_0_0_0_2/roundingadder/n151_o[0] ) );
  DFFX1 \fmul_0_0_0_0_3/roundingadder/n155_q_reg[0]  ( .D(
        \fmul_0_0_0_0_3/sigprodext [6]), .CLK(clk), .Q(
        \fmul_0_0_0_0_3/roundingadder/x_1_d1 [0]) );
  DFFX1 \fmul_0_0_0_0_3/roundingadder/n155_q_reg[1]  ( .D(
        \fmul_0_0_0_0_3/sigprodext [7]), .CLK(clk), .Q(
        \fmul_0_0_0_0_3/roundingadder/x_1_d1 [1]) );
  DFFX1 \fmul_0_0_0_0_3/roundingadder/n155_q_reg[2]  ( .D(
        \fmul_0_0_0_0_3/sigprodext [8]), .CLK(clk), .Q(
        \fmul_0_0_0_0_3/roundingadder/x_1_d1 [2]) );
  DFFX1 \fmul_0_0_0_0_3/roundingadder/n155_q_reg[3]  ( .D(
        \fmul_0_0_0_0_3/sigprodext [9]), .CLK(clk), .Q(
        \fmul_0_0_0_0_3/roundingadder/x_1_d1 [3]) );
  DFFX1 \fmul_0_0_0_0_3/roundingadder/n155_q_reg[4]  ( .D(
        \fmul_0_0_0_0_3/exppostnorm [0]), .CLK(clk), .Q(
        \fmul_0_0_0_0_3/roundingadder/x_1_d1 [4]) );
  DFFX1 \fmul_0_0_0_0_3/roundingadder/n155_q_reg[5]  ( .D(
        \fmul_0_0_0_0_3/exppostnorm [1]), .CLK(clk), .Q(
        \fmul_0_0_0_0_3/roundingadder/x_1_d1 [5]) );
  DFFX1 \fmul_0_0_0_0_3/roundingadder/n155_q_reg[6]  ( .D(
        \fmul_0_0_0_0_3/exppostnorm [2]), .CLK(clk), .Q(
        \fmul_0_0_0_0_3/roundingadder/x_1_d1 [6]) );
  DFFX1 \fmul_0_0_0_0_3/roundingadder/n155_q_reg[7]  ( .D(
        \fmul_0_0_0_0_3/exppostnorm [3]), .CLK(clk), .Q(
        \fmul_0_0_0_0_3/roundingadder/x_1_d1 [7]) );
  DFFX1 \fmul_0_0_0_0_3/roundingadder/n155_q_reg[8]  ( .D(
        \fmul_0_0_0_0_3/exppostnorm [4]), .CLK(clk), .Q(
        \fmul_0_0_0_0_3/roundingadder/x_1_d1 [8]) );
  DFFX1 \fmul_0_0_0_0_3/roundingadder/n155_q_reg[9]  ( .D(
        \fmul_0_0_0_0_3/exppostnorm [5]), .CLK(clk), .Q(
        \fmul_0_0_0_0_3/roundingadder/x_1_d1 [9]) );
  DFFX1 \fmul_0_0_0_0_3/roundingadder/n155_q_reg[10]  ( .D(n14134), .CLK(clk), 
        .Q(\fmul_0_0_0_0_3/roundingadder/x_1_d1 [10]) );
  DFFX1 \fmul_0_0_0_0_3/roundingadder/n154_q_reg  ( .D(\fmul_0_0_0_0_3/round ), 
        .CLK(clk), .Q(\fmul_0_0_0_0_3/roundingadder/n151_o[0] ) );
  DFFX1 \fadd_0_0_0_0_3_y_reg[0]  ( .D(n13111), .CLK(clk), .Q(n13638), .QN(
        n11677) );
  DFFX1 \fadd_0_0_0_0_3_y_reg[1]  ( .D(n13110), .CLK(clk), .Q(n13666), .QN(
        n11678) );
  DFFX1 \fadd_0_0_0_0_3_y_reg[2]  ( .D(n13109), .CLK(clk), .Q(n13687), .QN(
        n11679) );
  DFFX1 \fadd_0_0_0_0_3_y_reg[3]  ( .D(n13108), .CLK(clk), .Q(n13709), .QN(
        n11680) );
  DFFX1 \fadd_0_0_0_0_3_y_reg[4]  ( .D(n13107), .CLK(clk), .Q(n5766), .QN(
        n14568) );
  DFFX1 \fadd_0_0_0_0_3_y_reg[5]  ( .D(n13106), .CLK(clk), .Q(n5767), .QN(
        n14567) );
  DFFX1 \fadd_0_0_0_0_3_y_reg[6]  ( .D(n13105), .CLK(clk), .Q(n5768), .QN(
        n14566) );
  DFFX1 \fadd_0_0_0_0_3_y_reg[7]  ( .D(n13104), .CLK(clk), .Q(n5769), .QN(
        n14565) );
  DFFX1 \fadd_0_0_0_0_3_y_reg[8]  ( .D(n13103), .CLK(clk), .Q(n5770), .QN(
        n14564) );
  DFFX1 \fadd_0_0_0_0_3_y_reg[11]  ( .D(n13100), .CLK(clk), .Q(n13623), .QN(
        n12726) );
  DFFX1 \fadd_0_0_0_0_3_y_reg[10]  ( .D(n13101), .CLK(clk), .Q(n13890), .QN(
        n11687) );
  DFFX1 \fadd_0_0_0_0_3/n293_q_reg[0]  ( .D(\fadd_0_0_0_0_3/newy_10 ), .CLK(
        clk), .Q(\fadd_0_0_0_0_3/syncexnxy_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_3/n294_q_reg[0]  ( .D(\fadd_0_0_0_0_3/syncexnxy_d1 [0]), 
        .CLK(clk), .Q(n12329) );
  DFFX1 \p_val_107_reg[9]  ( .D(n12664), .CLK(clk), .Q(n13980) );
  DFFX1 \p_val_290_reg[9]  ( .D(n12663), .CLK(clk), .Q(n14105), .QN(n12324) );
  DFFX1 \fadd_0_0_0_0_2_y_reg[9]  ( .D(n13078), .CLK(clk), .QN(n11707) );
  DFFX1 \fadd_0_0_0_0_3_x_reg[9]  ( .D(n13090), .CLK(clk), .Q(n13580), .QN(
        n11697) );
  DFFX1 \fadd_0_0_0_0_3/n288_q_reg  ( .D(\fadd_0_0_0_0_3/newy_9 ), .CLK(clk), 
        .Q(\fadd_0_0_0_0_3/syncsigny_d1 ) );
  DFFX1 \fadd_0_0_0_0_3/n289_q_reg  ( .D(\fadd_0_0_0_0_3/syncsigny_d1 ), .CLK(
        clk), .QN(n12326) );
  DFFX1 \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[7]  ( .D(
        n12722), .CLK(clk), .Q(
        \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [7]) );
  DFFX1 \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[7]  ( .D(
        \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [7]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [7]) );
  DFFX1 \fadd_0_0_0_0_3/n284_q_reg  ( .D(n12722), .CLK(clk), .Q(
        \fadd_0_0_0_0_3/synceffsub_d1 ) );
  DFFX1 \fadd_0_0_0_0_3/n285_q_reg  ( .D(\fadd_0_0_0_0_3/synceffsub_d1 ), 
        .CLK(clk), .QN(n12320) );
  DFFX1 \fadd_0_0_0_0_3/n276_q_reg  ( .D(n12722), .CLK(clk), .Q(
        \fadd_0_0_0_0_3/effsub_d1 ) );
  DFFX1 \fadd_0_0_0_0_3/n277_q_reg  ( .D(\fadd_0_0_0_0_3/effsub_d1 ), .CLK(clk), .QN(n11518) );
  DFFX1 \p_val_107_reg[11]  ( .D(n12662), .CLK(clk), .Q(n13981) );
  DFFX1 \p_val_290_reg[11]  ( .D(n12661), .CLK(clk), .Q(n13840) );
  DFFX1 \fadd_0_0_0_0_2_y_reg[11]  ( .D(n13076), .CLK(clk), .Q(n13470), .QN(
        n12716) );
  DFFX1 \fadd_0_0_0_0_3_x_reg[11]  ( .D(n13088), .CLK(clk), .Q(n13510), .QN(
        n12724) );
  DFFX1 \fadd_0_0_0_0_3/n293_q_reg[3]  ( .D(\fadd_0_0_0_0_3/newx [11]), .CLK(
        clk), .Q(\fadd_0_0_0_0_3/syncexnxy_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_3/n294_q_reg[3]  ( .D(\fadd_0_0_0_0_3/syncexnxy_d1 [3]), 
        .CLK(clk), .Q(n13775), .QN(n12327) );
  DFFX1 \p_val_107_reg[10]  ( .D(n12660), .CLK(clk), .Q(n13982) );
  DFFX1 \p_val_290_reg[10]  ( .D(n12659), .CLK(clk), .Q(n13841) );
  DFFX1 \fadd_0_0_0_0_2_y_reg[10]  ( .D(n13077), .CLK(clk), .Q(n13589), .QN(
        n11708) );
  DFFX1 \fadd_0_0_0_0_3_x_reg[10]  ( .D(n13089), .CLK(clk), .Q(n13474), .QN(
        n12725) );
  DFFX1 \fadd_0_0_0_0_3/n286_q_reg[9]  ( .D(n14732), .CLK(clk), .Q(
        \fadd_0_0_0_0_3/syncx_d1 [9]) );
  DFFX1 \fadd_0_0_0_0_3/n287_q_reg[9]  ( .D(\fadd_0_0_0_0_3/syncx_d1 [9]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_3/syncx_d2 [9]) );
  DFFX1 \fadd_0_0_0_0_3/n286_q_reg[0]  ( .D(
        \add_0_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .CLK(clk), .Q(\fadd_0_0_0_0_3/syncx_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_3/n287_q_reg[0]  ( .D(\fadd_0_0_0_0_3/syncx_d1 [0]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_3/syncx_d2 [0]) );
  DFFX1 \p_val_107_reg[0]  ( .D(n12658), .CLK(clk), .Q(n13983) );
  DFFX1 \p_val_290_reg[0]  ( .D(n12657), .CLK(clk), .Q(n13870) );
  DFFX1 \fadd_0_0_0_0_2_y_reg[0]  ( .D(n13087), .CLK(clk), .Q(n13524), .QN(
        n11698) );
  DFFX1 \fadd_0_0_0_0_3_x_reg[0]  ( .D(n13099), .CLK(clk), .Q(n13518), .QN(
        n11688) );
  DFFX1 \fadd_0_0_0_0_3/rightshiftercomponent/n415_q_reg[2]  ( .D(n14736), 
        .CLK(clk), .QN(n11524) );
  DFFX1 \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/n432_q_reg[2]  ( .D(
        \add_0_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .CLK(clk), .Q(\fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/n433_q_reg[2]  ( .D(
        \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [2]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/x_d2 [2]) );
  DFFX1 \fadd_0_0_0_0_3/n293_q_reg[2]  ( .D(\fadd_0_0_0_0_3/newx [10]), .CLK(
        clk), .Q(\fadd_0_0_0_0_3/syncexnxy_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_3/n294_q_reg[2]  ( .D(\fadd_0_0_0_0_3/syncexnxy_d1 [2]), 
        .CLK(clk), .Q(n13731), .QN(n12325) );
  DFFX1 \fadd_0_0_0_0_3/n286_q_reg[1]  ( .D(
        \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ), .CLK(clk), .Q(\fadd_0_0_0_0_3/syncx_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_3/n287_q_reg[1]  ( .D(\fadd_0_0_0_0_3/syncx_d1 [1]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_3/syncx_d2 [1]) );
  DFFX1 \p_val_107_reg[1]  ( .D(n12656), .CLK(clk), .Q(n13984) );
  DFFX1 \p_val_290_reg[1]  ( .D(n12655), .CLK(clk), .Q(n13871) );
  DFFX1 \fadd_0_0_0_0_2_y_reg[1]  ( .D(n13086), .CLK(clk), .Q(n13535), .QN(
        n11699) );
  DFFX1 \fadd_0_0_0_0_3_x_reg[1]  ( .D(n13098), .CLK(clk), .Q(n13529), .QN(
        n11689) );
  DFFX1 \fadd_0_0_0_0_3/rightshiftercomponent/n415_q_reg[3]  ( .D(n14735), 
        .CLK(clk), .QN(n11525) );
  DFFX1 \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/n432_q_reg[3]  ( .D(
        \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ), .CLK(clk), .Q(\fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/n433_q_reg[3]  ( .D(
        \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [3]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/x_d2 [3]) );
  DFFX1 \fadd_0_0_0_0_3/n286_q_reg[2]  ( .D(
        \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ), .CLK(clk), .Q(\fadd_0_0_0_0_3/syncx_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_3/n287_q_reg[2]  ( .D(\fadd_0_0_0_0_3/syncx_d1 [2]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_3/syncx_d2 [2]) );
  DFFX1 \p_val_107_reg[2]  ( .D(n12654), .CLK(clk), .Q(n13985) );
  DFFX1 \p_val_290_reg[2]  ( .D(n12653), .CLK(clk), .Q(n13872) );
  DFFX1 \fadd_0_0_0_0_2_y_reg[2]  ( .D(n13085), .CLK(clk), .Q(n13560), .QN(
        n11700) );
  DFFX1 \fadd_0_0_0_0_3_x_reg[2]  ( .D(n13097), .CLK(clk), .Q(n13554), .QN(
        n11690) );
  DFFX1 \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/n432_q_reg[4]  ( .D(
        \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ), .CLK(clk), .Q(\fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/n433_q_reg[4]  ( .D(
        \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [4]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/x_d2 [4]) );
  DFFX1 \fadd_0_0_0_0_3/n286_q_reg[3]  ( .D(
        \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ), .CLK(clk), .Q(\fadd_0_0_0_0_3/syncx_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_3/n287_q_reg[3]  ( .D(\fadd_0_0_0_0_3/syncx_d1 [3]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_3/syncx_d2 [3]) );
  DFFX1 \p_val_107_reg[3]  ( .D(n12652), .CLK(clk), .Q(n13986) );
  DFFX1 \p_val_290_reg[3]  ( .D(n12651), .CLK(clk), .Q(n13873) );
  DFFX1 \fadd_0_0_0_0_2_y_reg[3]  ( .D(n13084), .CLK(clk), .Q(n13577), .QN(
        n11701) );
  DFFX1 \fadd_0_0_0_0_3_x_reg[3]  ( .D(n13096), .CLK(clk), .Q(n13571), .QN(
        n11691) );
  DFFX1 \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/n432_q_reg[5]  ( .D(
        \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ), .CLK(clk), .Q(\fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [5]) );
  DFFX1 \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/n433_q_reg[5]  ( .D(
        \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [5]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/x_d2 [5]) );
  DFFX1 \fadd_0_0_0_0_3/n275_q_reg[4]  ( .D(\fadd_0_0_0_0_3/newx [4]), .CLK(
        clk), .Q(\fadd_0_0_0_0_3/newx_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_3/n281_q_reg[0]  ( .D(\fadd_0_0_0_0_3/newx [4]), .CLK(
        clk), .Q(\fadd_0_0_0_0_3/exponentresultfar0_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_3/n282_q_reg[0]  ( .D(
        \fadd_0_0_0_0_3/exponentresultfar0_d1 [0]), .CLK(clk), .Q(
        \fadd_0_0_0_0_3/exponentresultfar0_d2 [0]) );
  DFFX1 \fadd_0_0_0_0_3/n286_q_reg[4]  ( .D(\fadd_0_0_0_0_3/newx [4]), .CLK(
        clk), .Q(\fadd_0_0_0_0_3/syncx_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_3/n287_q_reg[4]  ( .D(\fadd_0_0_0_0_3/syncx_d1 [4]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_3/syncx_d2 [4]) );
  DFFX1 \p_val_107_reg[4]  ( .D(n12650), .CLK(clk), .Q(n13987) );
  DFFX1 \p_val_290_reg[4]  ( .D(n12649), .CLK(clk), .Q(n13874) );
  DFFX1 \fadd_0_0_0_0_2_y_reg[4]  ( .D(n13083), .CLK(clk), .Q(n5838), .QN(
        n14557) );
  DFFX1 \fadd_0_0_0_0_3_x_reg[4]  ( .D(n13095), .CLK(clk), .Q(n5778), .QN(
        n14573) );
  DFFX1 \fadd_0_0_0_0_3/n275_q_reg[5]  ( .D(\fadd_0_0_0_0_3/newx [5]), .CLK(
        clk), .Q(\fadd_0_0_0_0_3/newx_d1 [5]) );
  DFFX1 \fadd_0_0_0_0_3/n281_q_reg[1]  ( .D(\fadd_0_0_0_0_3/newx [5]), .CLK(
        clk), .Q(\fadd_0_0_0_0_3/exponentresultfar0_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_3/n282_q_reg[1]  ( .D(
        \fadd_0_0_0_0_3/exponentresultfar0_d1 [1]), .CLK(clk), .Q(
        \fadd_0_0_0_0_3/exponentresultfar0_d2 [1]) );
  DFFX1 \fadd_0_0_0_0_3/n286_q_reg[5]  ( .D(\fadd_0_0_0_0_3/newx [5]), .CLK(
        clk), .Q(\fadd_0_0_0_0_3/syncx_d1 [5]) );
  DFFX1 \fadd_0_0_0_0_3/n287_q_reg[5]  ( .D(\fadd_0_0_0_0_3/syncx_d1 [5]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_3/syncx_d2 [5]) );
  DFFX1 \p_val_107_reg[5]  ( .D(n12648), .CLK(clk), .Q(n13988) );
  DFFX1 \p_val_290_reg[5]  ( .D(n12647), .CLK(clk), .Q(n13875) );
  DFFX1 \fadd_0_0_0_0_2_y_reg[5]  ( .D(n13082), .CLK(clk), .Q(n5839), .QN(
        n14556) );
  DFFX1 \fadd_0_0_0_0_3_x_reg[5]  ( .D(n13094), .CLK(clk), .Q(n5779), .QN(
        n14572) );
  DFFX1 \fadd_0_0_0_0_3/n275_q_reg[6]  ( .D(\fadd_0_0_0_0_3/newx [6]), .CLK(
        clk), .Q(\fadd_0_0_0_0_3/newx_d1 [6]) );
  DFFX1 \fadd_0_0_0_0_3/n281_q_reg[2]  ( .D(\fadd_0_0_0_0_3/newx [6]), .CLK(
        clk), .Q(\fadd_0_0_0_0_3/exponentresultfar0_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_3/n282_q_reg[2]  ( .D(
        \fadd_0_0_0_0_3/exponentresultfar0_d1 [2]), .CLK(clk), .Q(
        \fadd_0_0_0_0_3/exponentresultfar0_d2 [2]) );
  DFFX1 \fadd_0_0_0_0_3/n286_q_reg[6]  ( .D(\fadd_0_0_0_0_3/newx [6]), .CLK(
        clk), .Q(\fadd_0_0_0_0_3/syncx_d1 [6]) );
  DFFX1 \fadd_0_0_0_0_3/n287_q_reg[6]  ( .D(\fadd_0_0_0_0_3/syncx_d1 [6]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_3/syncx_d2 [6]) );
  DFFX1 \p_val_107_reg[6]  ( .D(n12646), .CLK(clk), .Q(n13989) );
  DFFX1 \p_val_290_reg[6]  ( .D(n12645), .CLK(clk), .Q(n13876) );
  DFFX1 \fadd_0_0_0_0_2_y_reg[6]  ( .D(n13081), .CLK(clk), .Q(n5840), .QN(
        n14555) );
  DFFX1 \fadd_0_0_0_0_3_x_reg[6]  ( .D(n13093), .CLK(clk), .Q(n5780), .QN(
        n14571) );
  DFFX1 \fadd_0_0_0_0_3/n275_q_reg[7]  ( .D(\fadd_0_0_0_0_3/newx [7]), .CLK(
        clk), .Q(\fadd_0_0_0_0_3/newx_d1 [7]) );
  DFFX1 \fadd_0_0_0_0_3/n281_q_reg[3]  ( .D(\fadd_0_0_0_0_3/newx [7]), .CLK(
        clk), .Q(\fadd_0_0_0_0_3/exponentresultfar0_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_3/n282_q_reg[3]  ( .D(
        \fadd_0_0_0_0_3/exponentresultfar0_d1 [3]), .CLK(clk), .Q(
        \fadd_0_0_0_0_3/exponentresultfar0_d2 [3]) );
  DFFX1 \fadd_0_0_0_0_3/n286_q_reg[7]  ( .D(\fadd_0_0_0_0_3/newx [7]), .CLK(
        clk), .Q(\fadd_0_0_0_0_3/syncx_d1 [7]) );
  DFFX1 \fadd_0_0_0_0_3/n287_q_reg[7]  ( .D(\fadd_0_0_0_0_3/syncx_d1 [7]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_3/syncx_d2 [7]) );
  DFFX1 \p_val_107_reg[7]  ( .D(n12644), .CLK(clk), .Q(n13990) );
  DFFX1 \p_val_290_reg[7]  ( .D(n12643), .CLK(clk), .Q(n13877) );
  DFFX1 \fadd_0_0_0_0_2_y_reg[7]  ( .D(n13080), .CLK(clk), .Q(n5841), .QN(
        n14554) );
  DFFX1 \fadd_0_0_0_0_3_x_reg[7]  ( .D(n13092), .CLK(clk), .Q(n5781), .QN(
        n14570) );
  DFFX1 \fadd_0_0_0_0_3/n275_q_reg[8]  ( .D(\fadd_0_0_0_0_3/newx [8]), .CLK(
        clk), .Q(\fadd_0_0_0_0_3/newx_d1 [8]) );
  DFFX1 \fadd_0_0_0_0_3/n280_q_reg[0]  ( .D(
        \fadd_0_0_0_0_3/exponentresultclose [0]), .CLK(clk), .Q(
        \fadd_0_0_0_0_3/exponentresultclose_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_3/n280_q_reg[1]  ( .D(
        \fadd_0_0_0_0_3/exponentresultclose [1]), .CLK(clk), .Q(
        \fadd_0_0_0_0_3/exponentresultclose_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_3/n280_q_reg[2]  ( .D(
        \fadd_0_0_0_0_3/exponentresultclose [2]), .CLK(clk), .Q(
        \fadd_0_0_0_0_3/exponentresultclose_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_3/n280_q_reg[3]  ( .D(
        \fadd_0_0_0_0_3/exponentresultclose [3]), .CLK(clk), .Q(
        \fadd_0_0_0_0_3/exponentresultclose_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_3/n280_q_reg[4]  ( .D(
        \fadd_0_0_0_0_3/exponentresultclose [4]), .CLK(clk), .Q(
        \fadd_0_0_0_0_3/exponentresultclose_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_3/n280_q_reg[6]  ( .D(n13662), .CLK(clk), .Q(
        \fadd_0_0_0_0_3/exponentresultclose_d1 [6]) );
  DFFX1 \fadd_0_0_0_0_3/n280_q_reg[5]  ( .D(n13662), .CLK(clk), .Q(
        \fadd_0_0_0_0_3/exponentresultclose_d1 [5]) );
  DFFX1 \fadd_0_0_0_0_3/n281_q_reg[4]  ( .D(\fadd_0_0_0_0_3/newx [8]), .CLK(
        clk), .Q(\fadd_0_0_0_0_3/exponentresultfar0_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_3/n282_q_reg[4]  ( .D(
        \fadd_0_0_0_0_3/exponentresultfar0_d1 [4]), .CLK(clk), .Q(
        \fadd_0_0_0_0_3/exponentresultfar0_d2 [4]) );
  DFFX1 \fadd_0_0_0_0_3/n286_q_reg[8]  ( .D(\fadd_0_0_0_0_3/newx [8]), .CLK(
        clk), .Q(\fadd_0_0_0_0_3/syncx_d1 [8]) );
  DFFX1 \fadd_0_0_0_0_3/n287_q_reg[8]  ( .D(\fadd_0_0_0_0_3/syncx_d1 [8]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_3/syncx_d2 [8]) );
  DFFX1 \p_val_107_reg[8]  ( .D(n12642), .CLK(clk), .Q(n13991) );
  DFFX1 \p_val_290_reg[8]  ( .D(n12641), .CLK(clk), .Q(n13878) );
  DFFX1 \fadd_0_0_0_0_2_y_reg[8]  ( .D(n13079), .CLK(clk), .Q(n5842), .QN(
        n14553) );
  DFFX1 \fadd_0_0_0_0_2/n275_q_reg[8]  ( .D(\fadd_0_0_0_0_2/newx [8]), .CLK(
        clk), .Q(\fadd_0_0_0_0_2/newx_d1 [8]) );
  DFFX1 \fadd_0_0_0_0_2/n281_q_reg[4]  ( .D(\fadd_0_0_0_0_2/newx [8]), .CLK(
        clk), .Q(\fadd_0_0_0_0_2/exponentresultfar0_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_2/n282_q_reg[4]  ( .D(
        \fadd_0_0_0_0_2/exponentresultfar0_d1 [4]), .CLK(clk), .Q(
        \fadd_0_0_0_0_2/exponentresultfar0_d2 [4]) );
  DFFX1 \fadd_0_0_0_0_2/n286_q_reg[8]  ( .D(\fadd_0_0_0_0_2/newx [8]), .CLK(
        clk), .Q(\fadd_0_0_0_0_2/syncx_d1 [8]) );
  DFFX1 \fadd_0_0_0_0_2/n287_q_reg[8]  ( .D(\fadd_0_0_0_0_2/syncx_d1 [8]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_2/syncx_d2 [8]) );
  DFFX1 \p_val_83_reg[8]  ( .D(n12640), .CLK(clk), .Q(n13917) );
  DFFX1 \p_val_289_reg[8]  ( .D(n12639), .CLK(clk), .Q(n13842) );
  DFFX1 \fadd_0_0_0_0_2_x_reg[8]  ( .D(n13067), .CLK(clk), .Q(n5854), .QN(
        n14562) );
  DFFX1 \fadd_0_0_0_0_2/rightshiftercomponent/n413_q_reg[0]  ( .D(n12711), 
        .CLK(clk), .Q(\fadd_0_0_0_0_2/rightshiftercomponent/ps_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_2/rightshiftercomponent/n414_q_reg[0]  ( .D(
        \fadd_0_0_0_0_2/rightshiftercomponent/ps_d1 [0]), .CLK(clk), .Q(
        \fadd_0_0_0_0_2/rightshiftercomponent/ps_d2[0] ) );
  DFFX1 \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[6]  ( .D(
        \fadd_0_0_0_0_2/fracyfarxorop [6]), .CLK(clk), .Q(
        \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [6]) );
  DFFX1 \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[6]  ( .D(
        \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [6]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [6]) );
  DFFX1 \p_val_83_reg[11]  ( .D(n12638), .CLK(clk), .Q(n13918) );
  DFFX1 \p_val_289_reg[11]  ( .D(n12637), .CLK(clk), .Q(n13843) );
  DFFX1 \fadd_0_0_0_0_2_x_reg[11]  ( .D(n13064), .CLK(clk), .Q(n13507), .QN(
        n12717) );
  DFFX1 \fadd_0_0_0_0_2/n293_q_reg[3]  ( .D(\fadd_0_0_0_0_2/newx [11]), .CLK(
        clk), .Q(\fadd_0_0_0_0_2/syncexnxy_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_2/n294_q_reg[3]  ( .D(\fadd_0_0_0_0_2/syncexnxy_d1 [3]), 
        .CLK(clk), .QN(n12297) );
  DFFX1 \p_val_83_reg[10]  ( .D(n12636), .CLK(clk), .Q(n13919) );
  DFFX1 \p_val_289_reg[10]  ( .D(n12635), .CLK(clk), .Q(n13844) );
  DFFX1 \fadd_0_0_0_0_2_x_reg[10]  ( .D(n13065), .CLK(clk), .Q(n13472), .QN(
        n12718) );
  DFFX1 \fadd_0_0_0_0_2/n293_q_reg[2]  ( .D(\fadd_0_0_0_0_2/newx [10]), .CLK(
        clk), .Q(\fadd_0_0_0_0_2/syncexnxy_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_2/n294_q_reg[2]  ( .D(\fadd_0_0_0_0_2/syncexnxy_d1 [2]), 
        .CLK(clk), .Q(n13727) );
  DFFX1 \fadd_0_0_0_0_2/n293_q_reg[0]  ( .D(\fadd_0_0_0_0_2/newy_10 ), .CLK(
        clk), .Q(\fadd_0_0_0_0_2/syncexnxy_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_2/n294_q_reg[0]  ( .D(\fadd_0_0_0_0_2/syncexnxy_d1 [0]), 
        .CLK(clk), .Q(n12299), .QN(n13738) );
  DFFX1 \fadd_0_0_0_0_2/n293_q_reg[1]  ( .D(\fadd_0_0_0_0_2/newy_11 ), .CLK(
        clk), .Q(\fadd_0_0_0_0_2/syncexnxy_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_2/n294_q_reg[1]  ( .D(\fadd_0_0_0_0_2/syncexnxy_d1 [1]), 
        .CLK(clk), .QN(n12298) );
  DFFX1 \p_val_83_reg[0]  ( .D(n12634), .CLK(clk), .Q(n13920) );
  DFFX1 \p_val_289_reg[0]  ( .D(n12633), .CLK(clk), .Q(n13845) );
  DFFX1 \fadd_0_0_0_0_2_x_reg[0]  ( .D(n13075), .CLK(clk), .Q(n13478), .QN(
        n11709) );
  DFFX1 \fadd_0_0_0_0_2/rightshiftercomponent/n415_q_reg[2]  ( .D(n14704), 
        .CLK(clk), .QN(n11511) );
  DFFX1 \fadd_0_0_0_0_2/n286_q_reg[0]  ( .D(
        \add_0_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .CLK(clk), .Q(\fadd_0_0_0_0_2/syncx_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_2/n287_q_reg[0]  ( .D(\fadd_0_0_0_0_2/syncx_d1 [0]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_2/syncx_d2 [0]) );
  DFFX1 \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/n432_q_reg[2]  ( .D(
        \add_0_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .CLK(clk), .Q(\fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/n433_q_reg[2]  ( .D(
        \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [2]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/x_d2 [2]) );
  DFFX1 \p_val_83_reg[1]  ( .D(n12632), .CLK(clk), .Q(n13921) );
  DFFX1 \p_val_289_reg[1]  ( .D(n12631), .CLK(clk), .Q(n13846) );
  DFFX1 \fadd_0_0_0_0_2_x_reg[1]  ( .D(n13074), .CLK(clk), .Q(n13480), .QN(
        n11710) );
  DFFX1 \fadd_0_0_0_0_2/rightshiftercomponent/n415_q_reg[3]  ( .D(n14703), 
        .CLK(clk), .QN(n11512) );
  DFFX1 \fadd_0_0_0_0_2/n286_q_reg[1]  ( .D(
        \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ), .CLK(clk), .Q(\fadd_0_0_0_0_2/syncx_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_2/n287_q_reg[1]  ( .D(\fadd_0_0_0_0_2/syncx_d1 [1]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_2/syncx_d2 [1]) );
  DFFX1 \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/n432_q_reg[3]  ( .D(
        \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ), .CLK(clk), .Q(\fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/n433_q_reg[3]  ( .D(
        \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [3]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/x_d2 [3]) );
  DFFX1 \p_val_83_reg[2]  ( .D(n12630), .CLK(clk), .Q(n13922) );
  DFFX1 \p_val_289_reg[2]  ( .D(n12629), .CLK(clk), .Q(n13847) );
  DFFX1 \fadd_0_0_0_0_2_x_reg[2]  ( .D(n13073), .CLK(clk), .Q(n13493), .QN(
        n11711) );
  DFFX1 \fadd_0_0_0_0_2/n286_q_reg[2]  ( .D(
        \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ), .CLK(clk), .Q(\fadd_0_0_0_0_2/syncx_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_2/n287_q_reg[2]  ( .D(\fadd_0_0_0_0_2/syncx_d1 [2]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_2/syncx_d2 [2]) );
  DFFX1 \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/n432_q_reg[4]  ( .D(
        \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ), .CLK(clk), .Q(\fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/n433_q_reg[4]  ( .D(
        \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [4]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/x_d2 [4]) );
  DFFX1 \p_val_83_reg[3]  ( .D(n12628), .CLK(clk), .Q(n13923) );
  DFFX1 \p_val_289_reg[3]  ( .D(n12627), .CLK(clk), .Q(n13848) );
  DFFX1 \fadd_0_0_0_0_2_x_reg[3]  ( .D(n13072), .CLK(clk), .Q(n13495), .QN(
        n11712) );
  DFFX1 \fadd_0_0_0_0_2/n286_q_reg[3]  ( .D(
        \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ), .CLK(clk), .Q(\fadd_0_0_0_0_2/syncx_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_2/n287_q_reg[3]  ( .D(\fadd_0_0_0_0_2/syncx_d1 [3]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_2/syncx_d2 [3]) );
  DFFX1 \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/n432_q_reg[5]  ( .D(
        \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ), .CLK(clk), .Q(\fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [5]) );
  DFFX1 \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/n433_q_reg[5]  ( .D(
        \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [5]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/x_d2 [5]) );
  DFFX1 \p_val_83_reg[4]  ( .D(n12626), .CLK(clk), .Q(n13924) );
  DFFX1 \p_val_289_reg[4]  ( .D(n12625), .CLK(clk), .Q(n13849) );
  DFFX1 \fadd_0_0_0_0_2_x_reg[4]  ( .D(n13071), .CLK(clk), .Q(n5850), .QN(
        n14561) );
  DFFX1 \fadd_0_0_0_0_2/n275_q_reg[4]  ( .D(\fadd_0_0_0_0_2/newx [4]), .CLK(
        clk), .Q(\fadd_0_0_0_0_2/newx_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_2/n281_q_reg[0]  ( .D(\fadd_0_0_0_0_2/newx [4]), .CLK(
        clk), .Q(\fadd_0_0_0_0_2/exponentresultfar0_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_2/n282_q_reg[0]  ( .D(
        \fadd_0_0_0_0_2/exponentresultfar0_d1 [0]), .CLK(clk), .Q(
        \fadd_0_0_0_0_2/exponentresultfar0_d2 [0]) );
  DFFX1 \fadd_0_0_0_0_2/n286_q_reg[4]  ( .D(\fadd_0_0_0_0_2/newx [4]), .CLK(
        clk), .Q(\fadd_0_0_0_0_2/syncx_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_2/n287_q_reg[4]  ( .D(\fadd_0_0_0_0_2/syncx_d1 [4]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_2/syncx_d2 [4]) );
  DFFX1 \p_val_83_reg[5]  ( .D(n12624), .CLK(clk), .Q(n13925) );
  DFFX1 \p_val_289_reg[5]  ( .D(n12623), .CLK(clk), .Q(n13850) );
  DFFX1 \fadd_0_0_0_0_2_x_reg[5]  ( .D(n13070), .CLK(clk), .Q(n5851), .QN(
        n14560) );
  DFFX1 \fadd_0_0_0_0_2/n275_q_reg[5]  ( .D(\fadd_0_0_0_0_2/newx [5]), .CLK(
        clk), .Q(\fadd_0_0_0_0_2/newx_d1 [5]) );
  DFFX1 \fadd_0_0_0_0_2/n281_q_reg[1]  ( .D(\fadd_0_0_0_0_2/newx [5]), .CLK(
        clk), .Q(\fadd_0_0_0_0_2/exponentresultfar0_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_2/n282_q_reg[1]  ( .D(
        \fadd_0_0_0_0_2/exponentresultfar0_d1 [1]), .CLK(clk), .Q(
        \fadd_0_0_0_0_2/exponentresultfar0_d2 [1]) );
  DFFX1 \fadd_0_0_0_0_2/n286_q_reg[5]  ( .D(\fadd_0_0_0_0_2/newx [5]), .CLK(
        clk), .Q(\fadd_0_0_0_0_2/syncx_d1 [5]) );
  DFFX1 \fadd_0_0_0_0_2/n287_q_reg[5]  ( .D(\fadd_0_0_0_0_2/syncx_d1 [5]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_2/syncx_d2 [5]) );
  DFFX1 \p_val_83_reg[6]  ( .D(n12622), .CLK(clk), .Q(n13926) );
  DFFX1 \p_val_289_reg[6]  ( .D(n12621), .CLK(clk), .Q(n13851) );
  DFFX1 \fadd_0_0_0_0_2_x_reg[6]  ( .D(n13069), .CLK(clk), .Q(n5852), .QN(
        n14559) );
  DFFX1 \fadd_0_0_0_0_2/n275_q_reg[6]  ( .D(\fadd_0_0_0_0_2/newx [6]), .CLK(
        clk), .Q(\fadd_0_0_0_0_2/newx_d1 [6]) );
  DFFX1 \fadd_0_0_0_0_2/n281_q_reg[2]  ( .D(\fadd_0_0_0_0_2/newx [6]), .CLK(
        clk), .Q(\fadd_0_0_0_0_2/exponentresultfar0_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_2/n282_q_reg[2]  ( .D(
        \fadd_0_0_0_0_2/exponentresultfar0_d1 [2]), .CLK(clk), .Q(
        \fadd_0_0_0_0_2/exponentresultfar0_d2 [2]) );
  DFFX1 \fadd_0_0_0_0_2/n286_q_reg[6]  ( .D(\fadd_0_0_0_0_2/newx [6]), .CLK(
        clk), .Q(\fadd_0_0_0_0_2/syncx_d1 [6]) );
  DFFX1 \fadd_0_0_0_0_2/n287_q_reg[6]  ( .D(\fadd_0_0_0_0_2/syncx_d1 [6]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_2/syncx_d2 [6]) );
  DFFX1 \p_val_83_reg[7]  ( .D(n12620), .CLK(clk), .Q(n13927) );
  DFFX1 \p_val_289_reg[7]  ( .D(n12619), .CLK(clk), .Q(n13852) );
  DFFX1 \fadd_0_0_0_0_2_x_reg[7]  ( .D(n13068), .CLK(clk), .Q(n5853), .QN(
        n14558) );
  DFFX1 \fadd_0_0_0_0_2/rightshiftercomponent/n413_q_reg[1]  ( .D(n14697), 
        .CLK(clk), .Q(\fadd_0_0_0_0_2/rightshiftercomponent/ps_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_2/rightshiftercomponent/n413_q_reg[2]  ( .D(n14694), 
        .CLK(clk), .Q(\fadd_0_0_0_0_2/rightshiftercomponent/ps_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_2/rightshiftercomponent/n416_q_reg[1]  ( .D(
        \fadd_0_0_0_0_2/rightshiftercomponent/level2[1] ), .CLK(clk), .QN(
        n11513) );
  DFFX1 \fadd_0_0_0_0_2/rightshiftercomponent/n416_q_reg[0]  ( .D(n12713), 
        .CLK(clk), .QN(n11514) );
  DFFX1 \fadd_0_0_0_0_2/rightshiftercomponent/n417_q_reg  ( .D(
        \fadd_0_0_0_0_2/rightshiftercomponent/n389_o ), .CLK(clk), .Q(n14946)
         );
  DFFX1 \fadd_0_0_0_0_2/rightshiftercomponent/n418_q_reg[0]  ( .D(n12712), 
        .CLK(clk), .Q(\fadd_0_0_0_0_2/rightshiftercomponent/level1_d1[0] ) );
  DFFX1 \fadd_0_0_0_0_2/rightshiftercomponent/n419_q_reg[0]  ( .D(
        \fadd_0_0_0_0_2/rightshiftercomponent/level1_d1[0] ), .CLK(clk), .Q(
        \fadd_0_0_0_0_2/rightshiftercomponent/level1_d2[0] ) );
  DFFX1 \fadd_0_0_0_0_2/n275_q_reg[7]  ( .D(\fadd_0_0_0_0_2/newx [7]), .CLK(
        clk), .Q(\fadd_0_0_0_0_2/newx_d1 [7]) );
  DFFX1 \fadd_0_0_0_0_2/n280_q_reg[0]  ( .D(
        \fadd_0_0_0_0_2/exponentresultclose [0]), .CLK(clk), .Q(
        \fadd_0_0_0_0_2/exponentresultclose_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_2/n280_q_reg[1]  ( .D(
        \fadd_0_0_0_0_2/exponentresultclose [1]), .CLK(clk), .Q(
        \fadd_0_0_0_0_2/exponentresultclose_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_2/n280_q_reg[2]  ( .D(
        \fadd_0_0_0_0_2/exponentresultclose [2]), .CLK(clk), .Q(
        \fadd_0_0_0_0_2/exponentresultclose_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_2/n280_q_reg[3]  ( .D(
        \fadd_0_0_0_0_2/exponentresultclose [3]), .CLK(clk), .Q(
        \fadd_0_0_0_0_2/exponentresultclose_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_2/n280_q_reg[4]  ( .D(
        \fadd_0_0_0_0_2/exponentresultclose [4]), .CLK(clk), .Q(
        \fadd_0_0_0_0_2/exponentresultclose_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_2/n280_q_reg[6]  ( .D(n13661), .CLK(clk), .Q(
        \fadd_0_0_0_0_2/exponentresultclose_d1 [6]) );
  DFFX1 \fadd_0_0_0_0_2/n280_q_reg[5]  ( .D(n13661), .CLK(clk), .Q(
        \fadd_0_0_0_0_2/exponentresultclose_d1 [5]) );
  DFFX1 \fadd_0_0_0_0_2/n281_q_reg[3]  ( .D(\fadd_0_0_0_0_2/newx [7]), .CLK(
        clk), .Q(\fadd_0_0_0_0_2/exponentresultfar0_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_2/n282_q_reg[3]  ( .D(
        \fadd_0_0_0_0_2/exponentresultfar0_d1 [3]), .CLK(clk), .Q(
        \fadd_0_0_0_0_2/exponentresultfar0_d2 [3]) );
  DFFX1 \fadd_0_0_0_0_2/n286_q_reg[7]  ( .D(\fadd_0_0_0_0_2/newx [7]), .CLK(
        clk), .Q(\fadd_0_0_0_0_2/syncx_d1 [7]) );
  DFFX1 \fadd_0_0_0_0_2/n287_q_reg[7]  ( .D(\fadd_0_0_0_0_2/syncx_d1 [7]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_2/syncx_d2 [7]) );
  DFFX1 \fadd_0_0_0_0_2/n278_q_reg  ( .D(n14693), .CLK(clk), .Q(
        \fadd_0_0_0_0_2/selectclosepath_d1 ), .QN(n11516) );
  DFFX1 \fadd_0_0_0_0_2/n283_q_reg  ( .D(\fadd_0_0_0_0_2/zerofromclose ), 
        .CLK(clk), .Q(\fadd_0_0_0_0_2/zerofromclose_d1 ) );
  DFFX1 \fadd_0_0_0_0_2/n290_q_reg  ( .D(\fadd_0_0_0_0_2/ressign ), .CLK(clk), 
        .Q(\fadd_0_0_0_0_2/syncressign_d1 ) );
  DFFX1 \fadd_0_0_0_0_2/n291_q_reg  ( .D(\fadd_0_0_0_0_2/syncressign_d1 ), 
        .CLK(clk), .QN(n12272) );
  DFFX1 \p_val_83_reg[9]  ( .D(n12618), .CLK(clk), .Q(n13928) );
  DFFX1 \p_val_289_reg[9]  ( .D(n12617), .CLK(clk), .QN(n12271) );
  DFFX1 \fadd_0_0_0_0_2_x_reg[9]  ( .D(n13066), .CLK(clk), .QN(n11718) );
  DFFX1 \fadd_0_0_0_0_2/n286_q_reg[9]  ( .D(n14700), .CLK(clk), .Q(
        \fadd_0_0_0_0_2/syncx_d1 [9]) );
  DFFX1 \fadd_0_0_0_0_2/n287_q_reg[9]  ( .D(\fadd_0_0_0_0_2/syncx_d1 [9]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_2/syncx_d2 [9]) );
  DFFX1 \fadd_0_0_0_0_2/n288_q_reg  ( .D(\fadd_0_0_0_0_2/newy_9 ), .CLK(clk), 
        .Q(\fadd_0_0_0_0_2/syncsigny_d1 ) );
  DFFX1 \fadd_0_0_0_0_2/n289_q_reg  ( .D(\fadd_0_0_0_0_2/syncsigny_d1 ), .CLK(
        clk), .Q(\fadd_0_0_0_0_2/syncsigny_d2 ) );
  DFFX1 \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[4]  ( .D(
        \fadd_0_0_0_0_2/fracyfarxorop [4]), .CLK(clk), .Q(
        \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[4]  ( .D(
        \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [4]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [4]) );
  DFFX1 \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[3]  ( .D(
        \fadd_0_0_0_0_2/fracyfarxorop [3]), .CLK(clk), .Q(
        \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[3]  ( .D(
        \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [3]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [3]) );
  DFFX1 \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[2]  ( .D(
        \fadd_0_0_0_0_2/fracyfarxorop [2]), .CLK(clk), .Q(
        \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[2]  ( .D(
        \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [2]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [2]) );
  DFFX1 \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[1]  ( .D(
        \fadd_0_0_0_0_2/fracyfarxorop [1]), .CLK(clk), .Q(
        \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[1]  ( .D(
        \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [1]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [1]) );
  DFFX1 \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[0]  ( .D(
        \fadd_0_0_0_0_2/fracyfarxorop [0]), .CLK(clk), .Q(
        \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[0]  ( .D(
        \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [0]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [0]) );
  DFFX1 \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[5]  ( .D(
        \fadd_0_0_0_0_2/fracyfarxorop [5]), .CLK(clk), .Q(
        \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [5]) );
  DFFX1 \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[5]  ( .D(
        \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [5]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [5]) );
  DFFX1 \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[7]  ( .D(
        n12714), .CLK(clk), .Q(
        \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [7]) );
  DFFX1 \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[7]  ( .D(
        \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [7]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [7]) );
  DFFX1 \fadd_0_0_0_0_2/n284_q_reg  ( .D(n12714), .CLK(clk), .Q(
        \fadd_0_0_0_0_2/synceffsub_d1 ) );
  DFFX1 \fadd_0_0_0_0_2/n285_q_reg  ( .D(\fadd_0_0_0_0_2/synceffsub_d1 ), 
        .CLK(clk), .QN(n12291) );
  DFFX1 \fadd_0_0_0_0_2/n276_q_reg  ( .D(n12714), .CLK(clk), .Q(
        \fadd_0_0_0_0_2/effsub_d1 ) );
  DFFX1 \fadd_0_0_0_0_2/n277_q_reg  ( .D(\fadd_0_0_0_0_2/effsub_d1 ), .CLK(clk), .QN(n11505) );
  DFFX1 \fadd_0_0_0_0_3_x_reg[8]  ( .D(n13091), .CLK(clk), .Q(n5782), .QN(
        n14569) );
  DFFX1 \fadd_0_0_0_0_3/rightshiftercomponent/n413_q_reg[2]  ( .D(n14726), 
        .CLK(clk), .Q(\fadd_0_0_0_0_3/rightshiftercomponent/ps_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_3/rightshiftercomponent/n416_q_reg[1]  ( .D(
        \fadd_0_0_0_0_3/rightshiftercomponent/level2[1] ), .CLK(clk), .QN(
        n11526) );
  DFFX1 \fadd_0_0_0_0_3/rightshiftercomponent/n416_q_reg[0]  ( .D(n12721), 
        .CLK(clk), .QN(n11527) );
  DFFX1 \fadd_0_0_0_0_3/rightshiftercomponent/n413_q_reg[1]  ( .D(n14729), 
        .CLK(clk), .Q(\fadd_0_0_0_0_3/rightshiftercomponent/ps_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_3/rightshiftercomponent/n417_q_reg  ( .D(
        \fadd_0_0_0_0_3/rightshiftercomponent/n389_o ), .CLK(clk), .Q(n14947)
         );
  DFFX1 \fadd_0_0_0_0_3/rightshiftercomponent/n418_q_reg[0]  ( .D(n12720), 
        .CLK(clk), .Q(\fadd_0_0_0_0_3/rightshiftercomponent/level1_d1[0] ) );
  DFFX1 \fadd_0_0_0_0_3/rightshiftercomponent/n419_q_reg[0]  ( .D(
        \fadd_0_0_0_0_3/rightshiftercomponent/level1_d1[0] ), .CLK(clk), .Q(
        \fadd_0_0_0_0_3/rightshiftercomponent/level1_d2[0] ) );
  DFFX1 \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[5]  ( .D(
        \fadd_0_0_0_0_3/fracyfarxorop [5]), .CLK(clk), .Q(
        \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [5]) );
  DFFX1 \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[5]  ( .D(
        \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [5]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [5]) );
  DFFX1 \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[3]  ( .D(
        \fadd_0_0_0_0_3/fracyfarxorop [3]), .CLK(clk), .Q(
        \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[3]  ( .D(
        \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [3]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [3]) );
  DFFX1 \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[2]  ( .D(
        \fadd_0_0_0_0_3/fracyfarxorop [2]), .CLK(clk), .Q(
        \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[2]  ( .D(
        \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [2]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [2]) );
  DFFX1 \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[1]  ( .D(
        \fadd_0_0_0_0_3/fracyfarxorop [1]), .CLK(clk), .Q(
        \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[1]  ( .D(
        \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [1]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [1]) );
  DFFX1 \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[0]  ( .D(
        \fadd_0_0_0_0_3/fracyfarxorop [0]), .CLK(clk), .Q(
        \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[0]  ( .D(
        \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [0]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [0]) );
  DFFX1 \fadd_0_0_0_0_3/rightshiftercomponent/n413_q_reg[0]  ( .D(n12719), 
        .CLK(clk), .Q(\fadd_0_0_0_0_3/rightshiftercomponent/ps_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_3/rightshiftercomponent/n414_q_reg[0]  ( .D(
        \fadd_0_0_0_0_3/rightshiftercomponent/ps_d1 [0]), .CLK(clk), .Q(
        \fadd_0_0_0_0_3/rightshiftercomponent/ps_d2[0] ) );
  DFFX1 \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[4]  ( .D(
        \fadd_0_0_0_0_3/fracyfarxorop [4]), .CLK(clk), .Q(
        \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[4]  ( .D(
        \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [4]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [4]) );
  DFFX1 \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[6]  ( .D(
        \fadd_0_0_0_0_3/fracyfarxorop [6]), .CLK(clk), .Q(
        \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [6]) );
  DFFX1 \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[6]  ( .D(
        \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [6]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [6]) );
  DFFX1 \fadd_0_0_0_0_3/n293_q_reg[1]  ( .D(\fadd_0_0_0_0_3/newy_11 ), .CLK(
        clk), .Q(\fadd_0_0_0_0_3/syncexnxy_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_3/n294_q_reg[1]  ( .D(\fadd_0_0_0_0_3/syncexnxy_d1 [1]), 
        .CLK(clk), .Q(n13740), .QN(n12328) );
  DFFX1 \fadd_0_0_0_0_3/n278_q_reg  ( .D(n14725), .CLK(clk), .Q(
        \fadd_0_0_0_0_3/selectclosepath_d1 ), .QN(n11529) );
  DFFX1 \fadd_0_0_0_0_3/n283_q_reg  ( .D(\fadd_0_0_0_0_3/zerofromclose ), 
        .CLK(clk), .Q(\fadd_0_0_0_0_3/zerofromclose_d1 ) );
  DFFX1 \fadd_0_0_0_0_3/n290_q_reg  ( .D(\fadd_0_0_0_0_3/ressign ), .CLK(clk), 
        .Q(\fadd_0_0_0_0_3/syncressign_d1 ) );
  DFFX1 \fadd_0_0_0_0_3/n291_q_reg  ( .D(\fadd_0_0_0_0_3/syncressign_d1 ), 
        .CLK(clk), .QN(n12330) );
  DFFX1 \fmul_0_0_0_0_4/roundingadder/n155_q_reg[0]  ( .D(
        \fmul_0_0_0_0_4/sigprodext [6]), .CLK(clk), .Q(
        \fmul_0_0_0_0_4/roundingadder/x_1_d1 [0]) );
  DFFX1 \fmul_0_0_0_0_4/roundingadder/n155_q_reg[1]  ( .D(
        \fmul_0_0_0_0_4/sigprodext [7]), .CLK(clk), .Q(
        \fmul_0_0_0_0_4/roundingadder/x_1_d1 [1]) );
  DFFX1 \fmul_0_0_0_0_4/roundingadder/n155_q_reg[2]  ( .D(
        \fmul_0_0_0_0_4/sigprodext [8]), .CLK(clk), .Q(
        \fmul_0_0_0_0_4/roundingadder/x_1_d1 [2]) );
  DFFX1 \fmul_0_0_0_0_4/roundingadder/n155_q_reg[3]  ( .D(
        \fmul_0_0_0_0_4/sigprodext [9]), .CLK(clk), .Q(
        \fmul_0_0_0_0_4/roundingadder/x_1_d1 [3]) );
  DFFX1 \fmul_0_0_0_0_4/roundingadder/n155_q_reg[4]  ( .D(
        \fmul_0_0_0_0_4/exppostnorm [0]), .CLK(clk), .Q(
        \fmul_0_0_0_0_4/roundingadder/x_1_d1 [4]) );
  DFFX1 \fmul_0_0_0_0_4/roundingadder/n155_q_reg[5]  ( .D(
        \fmul_0_0_0_0_4/exppostnorm [1]), .CLK(clk), .Q(
        \fmul_0_0_0_0_4/roundingadder/x_1_d1 [5]) );
  DFFX1 \fmul_0_0_0_0_4/roundingadder/n155_q_reg[6]  ( .D(
        \fmul_0_0_0_0_4/exppostnorm [2]), .CLK(clk), .Q(
        \fmul_0_0_0_0_4/roundingadder/x_1_d1 [6]) );
  DFFX1 \fmul_0_0_0_0_4/roundingadder/n155_q_reg[7]  ( .D(
        \fmul_0_0_0_0_4/exppostnorm [3]), .CLK(clk), .Q(
        \fmul_0_0_0_0_4/roundingadder/x_1_d1 [7]) );
  DFFX1 \fmul_0_0_0_0_4/roundingadder/n155_q_reg[8]  ( .D(
        \fmul_0_0_0_0_4/exppostnorm [4]), .CLK(clk), .Q(
        \fmul_0_0_0_0_4/roundingadder/x_1_d1 [8]) );
  DFFX1 \fmul_0_0_0_0_4/roundingadder/n155_q_reg[9]  ( .D(
        \fmul_0_0_0_0_4/exppostnorm [5]), .CLK(clk), .Q(
        \fmul_0_0_0_0_4/roundingadder/x_1_d1 [9]) );
  DFFX1 \fmul_0_0_0_0_4/roundingadder/n155_q_reg[10]  ( .D(n14133), .CLK(clk), 
        .Q(\fmul_0_0_0_0_4/roundingadder/x_1_d1 [10]) );
  DFFX1 \fmul_0_0_0_0_4/roundingadder/n154_q_reg  ( .D(\fmul_0_0_0_0_4/round ), 
        .CLK(clk), .Q(\fmul_0_0_0_0_4/roundingadder/n151_o[0] ) );
  DFFX1 \fmul_0_0_0_0_5/roundingadder/n155_q_reg[0]  ( .D(
        \fmul_0_0_0_0_5/sigprodext [6]), .CLK(clk), .Q(
        \fmul_0_0_0_0_5/roundingadder/x_1_d1 [0]) );
  DFFX1 \fmul_0_0_0_0_5/roundingadder/n155_q_reg[1]  ( .D(
        \fmul_0_0_0_0_5/sigprodext [7]), .CLK(clk), .Q(
        \fmul_0_0_0_0_5/roundingadder/x_1_d1 [1]) );
  DFFX1 \fmul_0_0_0_0_5/roundingadder/n155_q_reg[2]  ( .D(
        \fmul_0_0_0_0_5/sigprodext [8]), .CLK(clk), .Q(
        \fmul_0_0_0_0_5/roundingadder/x_1_d1 [2]) );
  DFFX1 \fmul_0_0_0_0_5/roundingadder/n155_q_reg[3]  ( .D(
        \fmul_0_0_0_0_5/sigprodext [9]), .CLK(clk), .Q(
        \fmul_0_0_0_0_5/roundingadder/x_1_d1 [3]) );
  DFFX1 \fmul_0_0_0_0_5/roundingadder/n155_q_reg[4]  ( .D(
        \fmul_0_0_0_0_5/exppostnorm [0]), .CLK(clk), .Q(
        \fmul_0_0_0_0_5/roundingadder/x_1_d1 [4]) );
  DFFX1 \fmul_0_0_0_0_5/roundingadder/n155_q_reg[5]  ( .D(
        \fmul_0_0_0_0_5/exppostnorm [1]), .CLK(clk), .Q(
        \fmul_0_0_0_0_5/roundingadder/x_1_d1 [5]) );
  DFFX1 \fmul_0_0_0_0_5/roundingadder/n155_q_reg[6]  ( .D(
        \fmul_0_0_0_0_5/exppostnorm [2]), .CLK(clk), .Q(
        \fmul_0_0_0_0_5/roundingadder/x_1_d1 [6]) );
  DFFX1 \fmul_0_0_0_0_5/roundingadder/n155_q_reg[7]  ( .D(
        \fmul_0_0_0_0_5/exppostnorm [3]), .CLK(clk), .Q(
        \fmul_0_0_0_0_5/roundingadder/x_1_d1 [7]) );
  DFFX1 \fmul_0_0_0_0_5/roundingadder/n155_q_reg[8]  ( .D(
        \fmul_0_0_0_0_5/exppostnorm [4]), .CLK(clk), .Q(
        \fmul_0_0_0_0_5/roundingadder/x_1_d1 [8]) );
  DFFX1 \fmul_0_0_0_0_5/roundingadder/n155_q_reg[9]  ( .D(
        \fmul_0_0_0_0_5/exppostnorm [5]), .CLK(clk), .Q(
        \fmul_0_0_0_0_5/roundingadder/x_1_d1 [9]) );
  DFFX1 \fmul_0_0_0_0_5/roundingadder/n155_q_reg[10]  ( .D(n14132), .CLK(clk), 
        .Q(\fmul_0_0_0_0_5/roundingadder/x_1_d1 [10]) );
  DFFX1 \fmul_0_0_0_0_5/roundingadder/n154_q_reg  ( .D(\fmul_0_0_0_0_5/round ), 
        .CLK(clk), .Q(\fmul_0_0_0_0_5/roundingadder/n151_o[0] ) );
  DFFX1 \fadd_0_0_0_0_5_y_reg[0]  ( .D(n13063), .CLK(clk), .Q(n13639), .QN(
        n11719) );
  DFFX1 \fadd_0_0_0_0_5_y_reg[1]  ( .D(n13062), .CLK(clk), .Q(n13667), .QN(
        n11720) );
  DFFX1 \fadd_0_0_0_0_5_y_reg[2]  ( .D(n13061), .CLK(clk), .Q(n13688), .QN(
        n11721) );
  DFFX1 \fadd_0_0_0_0_5_y_reg[3]  ( .D(n13060), .CLK(clk), .Q(n13710), .QN(
        n11722) );
  DFFX1 \fadd_0_0_0_0_5_y_reg[4]  ( .D(n13059), .CLK(clk), .Q(n5622), .QN(
        n14590) );
  DFFX1 \fadd_0_0_0_0_5_y_reg[5]  ( .D(n13058), .CLK(clk), .Q(n5623), .QN(
        n14589) );
  DFFX1 \fadd_0_0_0_0_5_y_reg[6]  ( .D(n13057), .CLK(clk), .Q(n5624), .QN(
        n14588) );
  DFFX1 \fadd_0_0_0_0_5_y_reg[7]  ( .D(n13056), .CLK(clk), .Q(n5625), .QN(
        n14587) );
  DFFX1 \fadd_0_0_0_0_5_y_reg[8]  ( .D(n13055), .CLK(clk), .Q(n5626), .QN(
        n14586) );
  DFFX1 \fadd_0_0_0_0_5_y_reg[11]  ( .D(n13052), .CLK(clk), .Q(n13624), .QN(
        n12746) );
  DFFX1 \fadd_0_0_0_0_5_y_reg[10]  ( .D(n13053), .CLK(clk), .Q(n13891), .QN(
        n11729) );
  DFFX1 \fadd_0_0_0_0_5/n293_q_reg[0]  ( .D(\fadd_0_0_0_0_5/newy_10 ), .CLK(
        clk), .Q(\fadd_0_0_0_0_5/syncexnxy_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_5/n294_q_reg[0]  ( .D(\fadd_0_0_0_0_5/syncexnxy_d1 [0]), 
        .CLK(clk), .Q(n12269), .QN(n13743) );
  DFFX1 \p_val_155_reg[0]  ( .D(n12616), .CLK(clk), .Q(n13992) );
  DFFX1 \p_val_292_reg[0]  ( .D(n12615), .CLK(clk), .Q(n13802) );
  DFFX1 \fadd_0_0_0_0_5_x_reg[0]  ( .D(n13051), .CLK(clk), .Q(n13519), .QN(
        n11730) );
  DFFX1 \fadd_0_0_0_0_5/n286_q_reg[0]  ( .D(
        \add_0_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .CLK(clk), .Q(\fadd_0_0_0_0_5/syncx_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_5/n287_q_reg[0]  ( .D(\fadd_0_0_0_0_5/syncx_d1 [0]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_5/syncx_d2 [0]) );
  DFFX1 \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/n432_q_reg[2]  ( .D(
        \add_0_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .CLK(clk), .Q(\fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/n433_q_reg[2]  ( .D(
        \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [2]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/x_d2 [2]) );
  DFFX1 \p_val_155_reg[11]  ( .D(n12614), .CLK(clk), .Q(n13993) );
  DFFX1 \p_val_292_reg[11]  ( .D(n12613), .CLK(clk), .Q(n13791) );
  DFFX1 \fadd_0_0_0_0_5_x_reg[11]  ( .D(n13040), .CLK(clk), .Q(n13511), .QN(
        n12744) );
  DFFX1 \fadd_0_0_0_0_5/n293_q_reg[3]  ( .D(\fadd_0_0_0_0_5/newx [11]), .CLK(
        clk), .Q(\fadd_0_0_0_0_5/syncexnxy_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_5/n294_q_reg[3]  ( .D(\fadd_0_0_0_0_5/syncexnxy_d1 [3]), 
        .CLK(clk), .Q(n13772), .QN(n12267) );
  DFFX1 \p_val_155_reg[10]  ( .D(n12612), .CLK(clk), .Q(n13994) );
  DFFX1 \p_val_292_reg[10]  ( .D(n12611), .CLK(clk), .Q(n13792) );
  DFFX1 \fadd_0_0_0_0_5_x_reg[10]  ( .D(n13041), .CLK(clk), .Q(n13503), .QN(
        n12745) );
  DFFX1 \fadd_0_0_0_0_5/rightshiftercomponent/n415_q_reg[2]  ( .D(n14789), 
        .CLK(clk), .QN(n11550) );
  DFFX1 \fadd_0_0_0_0_5/n293_q_reg[2]  ( .D(\fadd_0_0_0_0_5/newx [10]), .CLK(
        clk), .Q(\fadd_0_0_0_0_5/syncexnxy_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_5/n294_q_reg[2]  ( .D(\fadd_0_0_0_0_5/syncexnxy_d1 [2]), 
        .CLK(clk), .Q(n13733) );
  DFFX1 \fadd_0_0_0_0_5/n286_q_reg[1]  ( .D(
        \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ), .CLK(clk), .Q(\fadd_0_0_0_0_5/syncx_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_5/n287_q_reg[1]  ( .D(\fadd_0_0_0_0_5/syncx_d1 [1]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_5/syncx_d2 [1]) );
  DFFX1 \p_val_155_reg[1]  ( .D(n12610), .CLK(clk), .Q(n13995) );
  DFFX1 \p_val_292_reg[1]  ( .D(n12609), .CLK(clk), .Q(n13803) );
  DFFX1 \fadd_0_0_0_0_5_x_reg[1]  ( .D(n13050), .CLK(clk), .Q(n13530), .QN(
        n11731) );
  DFFX1 \fadd_0_0_0_0_5/rightshiftercomponent/n415_q_reg[3]  ( .D(n14788), 
        .CLK(clk), .QN(n11551) );
  DFFX1 \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/n432_q_reg[3]  ( .D(
        \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ), .CLK(clk), .Q(\fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/n433_q_reg[3]  ( .D(
        \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [3]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/x_d2 [3]) );
  DFFX1 \fadd_0_0_0_0_5/n286_q_reg[2]  ( .D(
        \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ), .CLK(clk), .Q(\fadd_0_0_0_0_5/syncx_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_5/n287_q_reg[2]  ( .D(\fadd_0_0_0_0_5/syncx_d1 [2]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_5/syncx_d2 [2]) );
  DFFX1 \p_val_155_reg[2]  ( .D(n12608), .CLK(clk), .Q(n13996) );
  DFFX1 \p_val_292_reg[2]  ( .D(n12607), .CLK(clk), .Q(n13804) );
  DFFX1 \fadd_0_0_0_0_5_x_reg[2]  ( .D(n13049), .CLK(clk), .Q(n13555), .QN(
        n11732) );
  DFFX1 \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/n432_q_reg[4]  ( .D(
        \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ), .CLK(clk), .Q(\fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/n433_q_reg[4]  ( .D(
        \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [4]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/x_d2 [4]) );
  DFFX1 \fadd_0_0_0_0_5/n286_q_reg[3]  ( .D(
        \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ), .CLK(clk), .Q(\fadd_0_0_0_0_5/syncx_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_5/n287_q_reg[3]  ( .D(\fadd_0_0_0_0_5/syncx_d1 [3]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_5/syncx_d2 [3]) );
  DFFX1 \p_val_155_reg[3]  ( .D(n12606), .CLK(clk), .Q(n13997) );
  DFFX1 \p_val_292_reg[3]  ( .D(n12605), .CLK(clk), .Q(n13805) );
  DFFX1 \fadd_0_0_0_0_5_x_reg[3]  ( .D(n13048), .CLK(clk), .Q(n13572), .QN(
        n11733) );
  DFFX1 \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/n432_q_reg[5]  ( .D(
        \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ), .CLK(clk), .Q(\fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [5]) );
  DFFX1 \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/n433_q_reg[5]  ( .D(
        \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [5]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/x_d2 [5]) );
  DFFX1 \fadd_0_0_0_0_5/n275_q_reg[4]  ( .D(\fadd_0_0_0_0_5/newx [4]), .CLK(
        clk), .Q(\fadd_0_0_0_0_5/newx_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_5/n281_q_reg[0]  ( .D(\fadd_0_0_0_0_5/newx [4]), .CLK(
        clk), .Q(\fadd_0_0_0_0_5/exponentresultfar0_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_5/n282_q_reg[0]  ( .D(
        \fadd_0_0_0_0_5/exponentresultfar0_d1 [0]), .CLK(clk), .Q(
        \fadd_0_0_0_0_5/exponentresultfar0_d2 [0]) );
  DFFX1 \fadd_0_0_0_0_5/n286_q_reg[4]  ( .D(\fadd_0_0_0_0_5/newx [4]), .CLK(
        clk), .Q(\fadd_0_0_0_0_5/syncx_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_5/n287_q_reg[4]  ( .D(\fadd_0_0_0_0_5/syncx_d1 [4]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_5/syncx_d2 [4]) );
  DFFX1 \p_val_155_reg[4]  ( .D(n12604), .CLK(clk), .Q(n13998) );
  DFFX1 \p_val_292_reg[4]  ( .D(n12603), .CLK(clk), .Q(n13806) );
  DFFX1 \fadd_0_0_0_0_5_x_reg[4]  ( .D(n13047), .CLK(clk), .Q(n5634), .QN(
        n14595) );
  DFFX1 \fadd_0_0_0_0_5/n275_q_reg[5]  ( .D(\fadd_0_0_0_0_5/newx [5]), .CLK(
        clk), .Q(\fadd_0_0_0_0_5/newx_d1 [5]) );
  DFFX1 \fadd_0_0_0_0_5/n281_q_reg[1]  ( .D(\fadd_0_0_0_0_5/newx [5]), .CLK(
        clk), .Q(\fadd_0_0_0_0_5/exponentresultfar0_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_5/n282_q_reg[1]  ( .D(
        \fadd_0_0_0_0_5/exponentresultfar0_d1 [1]), .CLK(clk), .Q(
        \fadd_0_0_0_0_5/exponentresultfar0_d2 [1]) );
  DFFX1 \fadd_0_0_0_0_5/n286_q_reg[5]  ( .D(\fadd_0_0_0_0_5/newx [5]), .CLK(
        clk), .Q(\fadd_0_0_0_0_5/syncx_d1 [5]) );
  DFFX1 \fadd_0_0_0_0_5/n287_q_reg[5]  ( .D(\fadd_0_0_0_0_5/syncx_d1 [5]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_5/syncx_d2 [5]) );
  DFFX1 \p_val_155_reg[5]  ( .D(n12602), .CLK(clk), .Q(n13999) );
  DFFX1 \p_val_292_reg[5]  ( .D(n12601), .CLK(clk), .Q(n13807) );
  DFFX1 \fadd_0_0_0_0_5_x_reg[5]  ( .D(n13046), .CLK(clk), .Q(n5635), .QN(
        n14594) );
  DFFX1 \fadd_0_0_0_0_5/n275_q_reg[6]  ( .D(\fadd_0_0_0_0_5/newx [6]), .CLK(
        clk), .Q(\fadd_0_0_0_0_5/newx_d1 [6]) );
  DFFX1 \fadd_0_0_0_0_5/n281_q_reg[2]  ( .D(\fadd_0_0_0_0_5/newx [6]), .CLK(
        clk), .Q(\fadd_0_0_0_0_5/exponentresultfar0_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_5/n282_q_reg[2]  ( .D(
        \fadd_0_0_0_0_5/exponentresultfar0_d1 [2]), .CLK(clk), .Q(
        \fadd_0_0_0_0_5/exponentresultfar0_d2 [2]) );
  DFFX1 \fadd_0_0_0_0_5/n286_q_reg[6]  ( .D(\fadd_0_0_0_0_5/newx [6]), .CLK(
        clk), .Q(\fadd_0_0_0_0_5/syncx_d1 [6]) );
  DFFX1 \fadd_0_0_0_0_5/n287_q_reg[6]  ( .D(\fadd_0_0_0_0_5/syncx_d1 [6]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_5/syncx_d2 [6]) );
  DFFX1 \p_val_155_reg[6]  ( .D(n12600), .CLK(clk), .Q(n14000) );
  DFFX1 \p_val_292_reg[6]  ( .D(n12599), .CLK(clk), .Q(n13808) );
  DFFX1 \fadd_0_0_0_0_5_x_reg[6]  ( .D(n13045), .CLK(clk), .Q(n5636), .QN(
        n14593) );
  DFFX1 \fadd_0_0_0_0_5/n275_q_reg[7]  ( .D(\fadd_0_0_0_0_5/newx [7]), .CLK(
        clk), .Q(\fadd_0_0_0_0_5/newx_d1 [7]) );
  DFFX1 \fadd_0_0_0_0_5/n281_q_reg[3]  ( .D(\fadd_0_0_0_0_5/newx [7]), .CLK(
        clk), .Q(\fadd_0_0_0_0_5/exponentresultfar0_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_5/n282_q_reg[3]  ( .D(
        \fadd_0_0_0_0_5/exponentresultfar0_d1 [3]), .CLK(clk), .Q(
        \fadd_0_0_0_0_5/exponentresultfar0_d2 [3]) );
  DFFX1 \fadd_0_0_0_0_5/n286_q_reg[7]  ( .D(\fadd_0_0_0_0_5/newx [7]), .CLK(
        clk), .Q(\fadd_0_0_0_0_5/syncx_d1 [7]) );
  DFFX1 \fadd_0_0_0_0_5/n287_q_reg[7]  ( .D(\fadd_0_0_0_0_5/syncx_d1 [7]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_5/syncx_d2 [7]) );
  DFFX1 \p_val_155_reg[7]  ( .D(n12598), .CLK(clk), .Q(n14001) );
  DFFX1 \p_val_292_reg[7]  ( .D(n12597), .CLK(clk), .Q(n13809) );
  DFFX1 \fadd_0_0_0_0_5_x_reg[7]  ( .D(n13044), .CLK(clk), .Q(n5637), .QN(
        n14592) );
  DFFX1 \fadd_0_0_0_0_5/n275_q_reg[8]  ( .D(\fadd_0_0_0_0_5/newx [8]), .CLK(
        clk), .Q(\fadd_0_0_0_0_5/newx_d1 [8]) );
  DFFX1 \fadd_0_0_0_0_5/n280_q_reg[0]  ( .D(
        \fadd_0_0_0_0_5/exponentresultclose [0]), .CLK(clk), .Q(
        \fadd_0_0_0_0_5/exponentresultclose_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_5/n280_q_reg[1]  ( .D(
        \fadd_0_0_0_0_5/exponentresultclose [1]), .CLK(clk), .Q(
        \fadd_0_0_0_0_5/exponentresultclose_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_5/n280_q_reg[2]  ( .D(
        \fadd_0_0_0_0_5/exponentresultclose [2]), .CLK(clk), .Q(
        \fadd_0_0_0_0_5/exponentresultclose_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_5/n280_q_reg[3]  ( .D(
        \fadd_0_0_0_0_5/exponentresultclose [3]), .CLK(clk), .Q(
        \fadd_0_0_0_0_5/exponentresultclose_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_5/n280_q_reg[4]  ( .D(
        \fadd_0_0_0_0_5/exponentresultclose [4]), .CLK(clk), .Q(
        \fadd_0_0_0_0_5/exponentresultclose_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_5/n280_q_reg[6]  ( .D(n13660), .CLK(clk), .Q(
        \fadd_0_0_0_0_5/exponentresultclose_d1 [6]) );
  DFFX1 \fadd_0_0_0_0_5/n280_q_reg[5]  ( .D(n13660), .CLK(clk), .Q(
        \fadd_0_0_0_0_5/exponentresultclose_d1 [5]) );
  DFFX1 \fadd_0_0_0_0_5/n281_q_reg[4]  ( .D(\fadd_0_0_0_0_5/newx [8]), .CLK(
        clk), .Q(\fadd_0_0_0_0_5/exponentresultfar0_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_5/n282_q_reg[4]  ( .D(
        \fadd_0_0_0_0_5/exponentresultfar0_d1 [4]), .CLK(clk), .Q(
        \fadd_0_0_0_0_5/exponentresultfar0_d2 [4]) );
  DFFX1 \fadd_0_0_0_0_5/n286_q_reg[8]  ( .D(\fadd_0_0_0_0_5/newx [8]), .CLK(
        clk), .Q(\fadd_0_0_0_0_5/syncx_d1 [8]) );
  DFFX1 \fadd_0_0_0_0_5/n287_q_reg[8]  ( .D(\fadd_0_0_0_0_5/syncx_d1 [8]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_5/syncx_d2 [8]) );
  DFFX1 \p_val_155_reg[8]  ( .D(n12596), .CLK(clk), .Q(n14002) );
  DFFX1 \p_val_292_reg[8]  ( .D(n12595), .CLK(clk), .Q(n13810) );
  DFFX1 \fadd_0_0_0_0_5_x_reg[8]  ( .D(n13043), .CLK(clk), .Q(n5638), .QN(
        n14591) );
  DFFX1 \fadd_0_0_0_0_5/rightshiftercomponent/n413_q_reg[2]  ( .D(n14779), 
        .CLK(clk), .Q(\fadd_0_0_0_0_5/rightshiftercomponent/ps_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_5/rightshiftercomponent/n416_q_reg[1]  ( .D(
        \fadd_0_0_0_0_5/rightshiftercomponent/level2[1] ), .CLK(clk), .QN(
        n11552) );
  DFFX1 \fadd_0_0_0_0_5/rightshiftercomponent/n416_q_reg[0]  ( .D(n12741), 
        .CLK(clk), .QN(n11553) );
  DFFX1 \fadd_0_0_0_0_5/rightshiftercomponent/n413_q_reg[1]  ( .D(n14782), 
        .CLK(clk), .Q(\fadd_0_0_0_0_5/rightshiftercomponent/ps_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_5/rightshiftercomponent/n417_q_reg  ( .D(
        \fadd_0_0_0_0_5/rightshiftercomponent/n389_o ), .CLK(clk), .Q(n14949)
         );
  DFFX1 \fadd_0_0_0_0_5/rightshiftercomponent/n418_q_reg[0]  ( .D(n12740), 
        .CLK(clk), .Q(\fadd_0_0_0_0_5/rightshiftercomponent/level1_d1[0] ) );
  DFFX1 \fadd_0_0_0_0_5/rightshiftercomponent/n419_q_reg[0]  ( .D(
        \fadd_0_0_0_0_5/rightshiftercomponent/level1_d1[0] ), .CLK(clk), .Q(
        \fadd_0_0_0_0_5/rightshiftercomponent/level1_d2[0] ) );
  DFFX1 \fadd_0_0_0_0_5/rightshiftercomponent/n413_q_reg[0]  ( .D(n12739), 
        .CLK(clk), .Q(\fadd_0_0_0_0_5/rightshiftercomponent/ps_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_5/rightshiftercomponent/n414_q_reg[0]  ( .D(
        \fadd_0_0_0_0_5/rightshiftercomponent/ps_d1 [0]), .CLK(clk), .Q(
        \fadd_0_0_0_0_5/rightshiftercomponent/ps_d2[0] ) );
  DFFX1 \fadd_0_0_0_0_5/n293_q_reg[1]  ( .D(\fadd_0_0_0_0_5/newy_11 ), .CLK(
        clk), .Q(\fadd_0_0_0_0_5/syncexnxy_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_5/n294_q_reg[1]  ( .D(\fadd_0_0_0_0_5/syncexnxy_d1 [1]), 
        .CLK(clk), .QN(n12268) );
  DFFX1 \fadd_0_0_0_0_5/n278_q_reg  ( .D(n14778), .CLK(clk), .Q(
        \fadd_0_0_0_0_5/selectclosepath_d1 ), .QN(n11555) );
  DFFX1 \fadd_0_0_0_0_5/n283_q_reg  ( .D(\fadd_0_0_0_0_5/zerofromclose ), 
        .CLK(clk), .Q(\fadd_0_0_0_0_5/zerofromclose_d1 ) );
  DFFX1 \fadd_0_0_0_0_5/n290_q_reg  ( .D(\fadd_0_0_0_0_5/ressign ), .CLK(clk), 
        .Q(\fadd_0_0_0_0_5/syncressign_d1 ) );
  DFFX1 \fadd_0_0_0_0_5/n291_q_reg  ( .D(\fadd_0_0_0_0_5/syncressign_d1 ), 
        .CLK(clk), .QN(n12242) );
  DFFX1 \p_val_155_reg[9]  ( .D(n12594), .CLK(clk), .Q(n14003) );
  DFFX1 \p_val_292_reg[9]  ( .D(n12593), .CLK(clk), .Q(n13779) );
  DFFX1 \fadd_0_0_0_0_5_x_reg[9]  ( .D(n13042), .CLK(clk), .Q(n13581), .QN(
        n11739) );
  DFFX1 \fadd_0_0_0_0_5/n286_q_reg[9]  ( .D(n14785), .CLK(clk), .Q(
        \fadd_0_0_0_0_5/syncx_d1 [9]) );
  DFFX1 \fadd_0_0_0_0_5/n287_q_reg[9]  ( .D(\fadd_0_0_0_0_5/syncx_d1 [9]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_5/syncx_d2 [9]) );
  DFFX1 \fadd_0_0_0_0_5/n288_q_reg  ( .D(\fadd_0_0_0_0_5/newy_9 ), .CLK(clk), 
        .Q(\fadd_0_0_0_0_5/syncsigny_d1 ) );
  DFFX1 \fadd_0_0_0_0_5/n289_q_reg  ( .D(\fadd_0_0_0_0_5/syncsigny_d1 ), .CLK(
        clk), .Q(\fadd_0_0_0_0_5/syncsigny_d2 ) );
  DFFX1 \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[6]  ( .D(
        \fadd_0_0_0_0_5/fracyfarxorop [6]), .CLK(clk), .Q(
        \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [6]) );
  DFFX1 \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[6]  ( .D(
        \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [6]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [6]) );
  DFFX1 \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[4]  ( .D(
        \fadd_0_0_0_0_5/fracyfarxorop [4]), .CLK(clk), .Q(
        \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[4]  ( .D(
        \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [4]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [4]) );
  DFFX1 \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[3]  ( .D(
        \fadd_0_0_0_0_5/fracyfarxorop [3]), .CLK(clk), .Q(
        \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[3]  ( .D(
        \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [3]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [3]) );
  DFFX1 \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[2]  ( .D(
        \fadd_0_0_0_0_5/fracyfarxorop [2]), .CLK(clk), .Q(
        \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[2]  ( .D(
        \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [2]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [2]) );
  DFFX1 \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[1]  ( .D(
        \fadd_0_0_0_0_5/fracyfarxorop [1]), .CLK(clk), .Q(
        \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[1]  ( .D(
        \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [1]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [1]) );
  DFFX1 \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[0]  ( .D(
        \fadd_0_0_0_0_5/fracyfarxorop [0]), .CLK(clk), .Q(
        \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[0]  ( .D(
        \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [0]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [0]) );
  DFFX1 \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[5]  ( .D(
        \fadd_0_0_0_0_5/fracyfarxorop [5]), .CLK(clk), .Q(
        \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [5]) );
  DFFX1 \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[5]  ( .D(
        \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [5]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [5]) );
  DFFX1 \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[7]  ( .D(
        n12742), .CLK(clk), .Q(
        \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [7]) );
  DFFX1 \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[7]  ( .D(
        \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [7]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [7]) );
  DFFX1 \fadd_0_0_0_0_5/n284_q_reg  ( .D(n12742), .CLK(clk), .Q(
        \fadd_0_0_0_0_5/synceffsub_d1 ) );
  DFFX1 \fadd_0_0_0_0_5/n285_q_reg  ( .D(\fadd_0_0_0_0_5/synceffsub_d1 ), 
        .CLK(clk), .QN(n12261) );
  DFFX1 \fadd_0_0_0_0_5/n276_q_reg  ( .D(n12742), .CLK(clk), .Q(
        \fadd_0_0_0_0_5/effsub_d1 ) );
  DFFX1 \fadd_0_0_0_0_5/n277_q_reg  ( .D(\fadd_0_0_0_0_5/effsub_d1 ), .CLK(clk), .QN(n11544) );
  DFFX1 \fmul_0_0_0_0_6/roundingadder/n155_q_reg[0]  ( .D(
        \fmul_0_0_0_0_6/sigprodext [6]), .CLK(clk), .Q(
        \fmul_0_0_0_0_6/roundingadder/x_1_d1 [0]) );
  DFFX1 \fmul_0_0_0_0_6/roundingadder/n155_q_reg[1]  ( .D(
        \fmul_0_0_0_0_6/sigprodext [7]), .CLK(clk), .Q(
        \fmul_0_0_0_0_6/roundingadder/x_1_d1 [1]) );
  DFFX1 \fmul_0_0_0_0_6/roundingadder/n155_q_reg[2]  ( .D(
        \fmul_0_0_0_0_6/sigprodext [8]), .CLK(clk), .Q(
        \fmul_0_0_0_0_6/roundingadder/x_1_d1 [2]) );
  DFFX1 \fmul_0_0_0_0_6/roundingadder/n155_q_reg[3]  ( .D(
        \fmul_0_0_0_0_6/sigprodext [9]), .CLK(clk), .Q(
        \fmul_0_0_0_0_6/roundingadder/x_1_d1 [3]) );
  DFFX1 \fmul_0_0_0_0_6/roundingadder/n155_q_reg[4]  ( .D(
        \fmul_0_0_0_0_6/exppostnorm [0]), .CLK(clk), .Q(
        \fmul_0_0_0_0_6/roundingadder/x_1_d1 [4]) );
  DFFX1 \fmul_0_0_0_0_6/roundingadder/n155_q_reg[5]  ( .D(
        \fmul_0_0_0_0_6/exppostnorm [1]), .CLK(clk), .Q(
        \fmul_0_0_0_0_6/roundingadder/x_1_d1 [5]) );
  DFFX1 \fmul_0_0_0_0_6/roundingadder/n155_q_reg[6]  ( .D(
        \fmul_0_0_0_0_6/exppostnorm [2]), .CLK(clk), .Q(
        \fmul_0_0_0_0_6/roundingadder/x_1_d1 [6]) );
  DFFX1 \fmul_0_0_0_0_6/roundingadder/n155_q_reg[7]  ( .D(
        \fmul_0_0_0_0_6/exppostnorm [3]), .CLK(clk), .Q(
        \fmul_0_0_0_0_6/roundingadder/x_1_d1 [7]) );
  DFFX1 \fmul_0_0_0_0_6/roundingadder/n155_q_reg[8]  ( .D(
        \fmul_0_0_0_0_6/exppostnorm [4]), .CLK(clk), .Q(
        \fmul_0_0_0_0_6/roundingadder/x_1_d1 [8]) );
  DFFX1 \fmul_0_0_0_0_6/roundingadder/n155_q_reg[9]  ( .D(
        \fmul_0_0_0_0_6/exppostnorm [5]), .CLK(clk), .Q(
        \fmul_0_0_0_0_6/roundingadder/x_1_d1 [9]) );
  DFFX1 \fmul_0_0_0_0_6/roundingadder/n155_q_reg[10]  ( .D(n14131), .CLK(clk), 
        .Q(\fmul_0_0_0_0_6/roundingadder/x_1_d1 [10]) );
  DFFX1 \fmul_0_0_0_0_6/roundingadder/n154_q_reg  ( .D(\fmul_0_0_0_0_6/round ), 
        .CLK(clk), .Q(\fmul_0_0_0_0_6/roundingadder/n151_o[0] ) );
  DFFX1 \fmul_0_0_0_0_7/roundingadder/n155_q_reg[0]  ( .D(
        \fmul_0_0_0_0_7/sigprodext [6]), .CLK(clk), .Q(
        \fmul_0_0_0_0_7/roundingadder/x_1_d1 [0]) );
  DFFX1 \fmul_0_0_0_0_7/roundingadder/n155_q_reg[1]  ( .D(
        \fmul_0_0_0_0_7/sigprodext [7]), .CLK(clk), .Q(
        \fmul_0_0_0_0_7/roundingadder/x_1_d1 [1]) );
  DFFX1 \fmul_0_0_0_0_7/roundingadder/n155_q_reg[2]  ( .D(
        \fmul_0_0_0_0_7/sigprodext [8]), .CLK(clk), .Q(
        \fmul_0_0_0_0_7/roundingadder/x_1_d1 [2]) );
  DFFX1 \fmul_0_0_0_0_7/roundingadder/n155_q_reg[3]  ( .D(
        \fmul_0_0_0_0_7/sigprodext [9]), .CLK(clk), .Q(
        \fmul_0_0_0_0_7/roundingadder/x_1_d1 [3]) );
  DFFX1 \fmul_0_0_0_0_7/roundingadder/n155_q_reg[4]  ( .D(
        \fmul_0_0_0_0_7/exppostnorm [0]), .CLK(clk), .Q(
        \fmul_0_0_0_0_7/roundingadder/x_1_d1 [4]) );
  DFFX1 \fmul_0_0_0_0_7/roundingadder/n155_q_reg[5]  ( .D(
        \fmul_0_0_0_0_7/exppostnorm [1]), .CLK(clk), .Q(
        \fmul_0_0_0_0_7/roundingadder/x_1_d1 [5]) );
  DFFX1 \fmul_0_0_0_0_7/roundingadder/n155_q_reg[6]  ( .D(
        \fmul_0_0_0_0_7/exppostnorm [2]), .CLK(clk), .Q(
        \fmul_0_0_0_0_7/roundingadder/x_1_d1 [6]) );
  DFFX1 \fmul_0_0_0_0_7/roundingadder/n155_q_reg[7]  ( .D(
        \fmul_0_0_0_0_7/exppostnorm [3]), .CLK(clk), .Q(
        \fmul_0_0_0_0_7/roundingadder/x_1_d1 [7]) );
  DFFX1 \fmul_0_0_0_0_7/roundingadder/n155_q_reg[8]  ( .D(
        \fmul_0_0_0_0_7/exppostnorm [4]), .CLK(clk), .Q(
        \fmul_0_0_0_0_7/roundingadder/x_1_d1 [8]) );
  DFFX1 \fmul_0_0_0_0_7/roundingadder/n155_q_reg[9]  ( .D(
        \fmul_0_0_0_0_7/exppostnorm [5]), .CLK(clk), .Q(
        \fmul_0_0_0_0_7/roundingadder/x_1_d1 [9]) );
  DFFX1 \fmul_0_0_0_0_7/roundingadder/n155_q_reg[10]  ( .D(n14130), .CLK(clk), 
        .Q(\fmul_0_0_0_0_7/roundingadder/x_1_d1 [10]) );
  DFFX1 \fmul_0_0_0_0_7/roundingadder/n154_q_reg  ( .D(\fmul_0_0_0_0_7/round ), 
        .CLK(clk), .Q(\fmul_0_0_0_0_7/roundingadder/n151_o[0] ) );
  DFFX1 \fadd_0_0_0_0_7_y_reg[0]  ( .D(n13039), .CLK(clk), .Q(n13640), .QN(
        n11740) );
  DFFX1 \fadd_0_0_0_0_7_y_reg[1]  ( .D(n13038), .CLK(clk), .Q(n13668), .QN(
        n11741) );
  DFFX1 \fadd_0_0_0_0_7_y_reg[2]  ( .D(n13037), .CLK(clk), .Q(n13689), .QN(
        n11742) );
  DFFX1 \fadd_0_0_0_0_7_y_reg[3]  ( .D(n13036), .CLK(clk), .Q(n13711), .QN(
        n11743) );
  DFFX1 \fadd_0_0_0_0_7_y_reg[4]  ( .D(n13035), .CLK(clk), .Q(n5478), .QN(
        n14612) );
  DFFX1 \fadd_0_0_0_0_7_y_reg[5]  ( .D(n13034), .CLK(clk), .Q(n5479), .QN(
        n14611) );
  DFFX1 \fadd_0_0_0_0_7_y_reg[6]  ( .D(n13033), .CLK(clk), .Q(n5480), .QN(
        n14610) );
  DFFX1 \fadd_0_0_0_0_7_y_reg[7]  ( .D(n13032), .CLK(clk), .Q(n5481), .QN(
        n14609) );
  DFFX1 \fadd_0_0_0_0_7_y_reg[8]  ( .D(n13031), .CLK(clk), .Q(n5482), .QN(
        n14608) );
  DFFX1 \fadd_0_0_0_0_7_y_reg[11]  ( .D(n13028), .CLK(clk), .Q(n13625), .QN(
        n12766) );
  DFFX1 \fadd_0_0_0_0_7_y_reg[10]  ( .D(n13029), .CLK(clk), .Q(n13892), .QN(
        n11750) );
  DFFX1 \fadd_0_0_0_0_7/n293_q_reg[0]  ( .D(\fadd_0_0_0_0_7/newy_10 ), .CLK(
        clk), .Q(\fadd_0_0_0_0_7/syncexnxy_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_7/n294_q_reg[0]  ( .D(\fadd_0_0_0_0_7/syncexnxy_d1 [0]), 
        .CLK(clk), .Q(n12239), .QN(n13744) );
  DFFX1 \p_val_203_reg[0]  ( .D(n12592), .CLK(clk), .Q(n14004) );
  DFFX1 \p_val_294_reg[0]  ( .D(n12591), .CLK(clk), .Q(n13853) );
  DFFX1 \fadd_0_0_0_0_6_y_reg[0]  ( .D(n13015), .CLK(clk), .Q(n13525), .QN(
        n11761) );
  DFFX1 \fadd_0_0_0_0_7_x_reg[0]  ( .D(n13027), .CLK(clk), .Q(n13520), .QN(
        n11751) );
  DFFX1 \fadd_0_0_0_0_7/n286_q_reg[0]  ( .D(
        \add_0_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .CLK(clk), .Q(\fadd_0_0_0_0_7/syncx_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_7/n287_q_reg[0]  ( .D(\fadd_0_0_0_0_7/syncx_d1 [0]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_7/syncx_d2 [0]) );
  DFFX1 \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/n432_q_reg[2]  ( .D(
        \add_0_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .CLK(clk), .Q(\fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/n433_q_reg[2]  ( .D(
        \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [2]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/x_d2 [2]) );
  DFFX1 \p_val_203_reg[11]  ( .D(n12590), .CLK(clk), .Q(n14005) );
  DFFX1 \p_val_294_reg[11]  ( .D(n12589), .CLK(clk), .Q(n13854) );
  DFFX1 \fadd_0_0_0_0_6_y_reg[11]  ( .D(n13004), .CLK(clk), .Q(n13471), .QN(
        n12756) );
  DFFX1 \fadd_0_0_0_0_7_x_reg[11]  ( .D(n13016), .CLK(clk), .Q(n13512), .QN(
        n12764) );
  DFFX1 \fadd_0_0_0_0_7/n293_q_reg[3]  ( .D(\fadd_0_0_0_0_7/newx [11]), .CLK(
        clk), .Q(\fadd_0_0_0_0_7/syncexnxy_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_7/n294_q_reg[3]  ( .D(\fadd_0_0_0_0_7/syncexnxy_d1 [3]), 
        .CLK(clk), .Q(n13773), .QN(n12237) );
  DFFX1 \p_val_203_reg[10]  ( .D(n12588), .CLK(clk), .Q(n14006) );
  DFFX1 \p_val_294_reg[10]  ( .D(n12587), .CLK(clk), .Q(n13857) );
  DFFX1 \fadd_0_0_0_0_6_y_reg[10]  ( .D(n13005), .CLK(clk), .Q(n13590), .QN(
        n11771) );
  DFFX1 \fadd_0_0_0_0_7_x_reg[10]  ( .D(n13017), .CLK(clk), .Q(n13475), .QN(
        n12765) );
  DFFX1 \fadd_0_0_0_0_7/rightshiftercomponent/n415_q_reg[2]  ( .D(n14831), 
        .CLK(clk), .QN(n11576) );
  DFFX1 \fadd_0_0_0_0_7/n293_q_reg[2]  ( .D(\fadd_0_0_0_0_7/newx [10]), .CLK(
        clk), .Q(\fadd_0_0_0_0_7/syncexnxy_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_7/n294_q_reg[2]  ( .D(\fadd_0_0_0_0_7/syncexnxy_d1 [2]), 
        .CLK(clk), .Q(n13734) );
  DFFX1 \fadd_0_0_0_0_7/n286_q_reg[1]  ( .D(
        \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ), .CLK(clk), .Q(\fadd_0_0_0_0_7/syncx_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_7/n287_q_reg[1]  ( .D(\fadd_0_0_0_0_7/syncx_d1 [1]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_7/syncx_d2 [1]) );
  DFFX1 \p_val_203_reg[1]  ( .D(n12586), .CLK(clk), .Q(n14007) );
  DFFX1 \p_val_294_reg[1]  ( .D(n12585), .CLK(clk), .Q(n13879) );
  DFFX1 \fadd_0_0_0_0_6_y_reg[1]  ( .D(n13014), .CLK(clk), .Q(n13536), .QN(
        n11762) );
  DFFX1 \fadd_0_0_0_0_7_x_reg[1]  ( .D(n13026), .CLK(clk), .Q(n13531), .QN(
        n11752) );
  DFFX1 \fadd_0_0_0_0_7/rightshiftercomponent/n415_q_reg[3]  ( .D(n14830), 
        .CLK(clk), .QN(n11577) );
  DFFX1 \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/n432_q_reg[3]  ( .D(
        \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ), .CLK(clk), .Q(\fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/n433_q_reg[3]  ( .D(
        \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [3]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/x_d2 [3]) );
  DFFX1 \fadd_0_0_0_0_7/n286_q_reg[2]  ( .D(
        \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ), .CLK(clk), .Q(\fadd_0_0_0_0_7/syncx_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_7/n287_q_reg[2]  ( .D(\fadd_0_0_0_0_7/syncx_d1 [2]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_7/syncx_d2 [2]) );
  DFFX1 \p_val_203_reg[2]  ( .D(n12584), .CLK(clk), .Q(n14008) );
  DFFX1 \p_val_294_reg[2]  ( .D(n12583), .CLK(clk), .Q(n13855) );
  DFFX1 \fadd_0_0_0_0_6_y_reg[2]  ( .D(n13013), .CLK(clk), .Q(n13561), .QN(
        n11763) );
  DFFX1 \fadd_0_0_0_0_7_x_reg[2]  ( .D(n13025), .CLK(clk), .Q(n13556), .QN(
        n11753) );
  DFFX1 \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/n432_q_reg[4]  ( .D(
        \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ), .CLK(clk), .Q(\fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/n433_q_reg[4]  ( .D(
        \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [4]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/x_d2 [4]) );
  DFFX1 \fadd_0_0_0_0_7/n286_q_reg[3]  ( .D(
        \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ), .CLK(clk), .Q(\fadd_0_0_0_0_7/syncx_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_7/n287_q_reg[3]  ( .D(\fadd_0_0_0_0_7/syncx_d1 [3]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_7/syncx_d2 [3]) );
  DFFX1 \p_val_203_reg[3]  ( .D(n12582), .CLK(clk), .Q(n14009) );
  DFFX1 \p_val_294_reg[3]  ( .D(n12581), .CLK(clk), .Q(n13880) );
  DFFX1 \fadd_0_0_0_0_6_y_reg[3]  ( .D(n13012), .CLK(clk), .Q(n13578), .QN(
        n11764) );
  DFFX1 \fadd_0_0_0_0_7_x_reg[3]  ( .D(n13024), .CLK(clk), .Q(n13573), .QN(
        n11754) );
  DFFX1 \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/n432_q_reg[5]  ( .D(
        \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ), .CLK(clk), .Q(\fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [5]) );
  DFFX1 \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/n433_q_reg[5]  ( .D(
        \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [5]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/x_d2 [5]) );
  DFFX1 \fadd_0_0_0_0_7/n275_q_reg[4]  ( .D(\fadd_0_0_0_0_7/newx [4]), .CLK(
        clk), .Q(\fadd_0_0_0_0_7/newx_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_7/n281_q_reg[0]  ( .D(\fadd_0_0_0_0_7/newx [4]), .CLK(
        clk), .Q(\fadd_0_0_0_0_7/exponentresultfar0_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_7/n282_q_reg[0]  ( .D(
        \fadd_0_0_0_0_7/exponentresultfar0_d1 [0]), .CLK(clk), .Q(
        \fadd_0_0_0_0_7/exponentresultfar0_d2 [0]) );
  DFFX1 \fadd_0_0_0_0_7/n286_q_reg[4]  ( .D(\fadd_0_0_0_0_7/newx [4]), .CLK(
        clk), .Q(\fadd_0_0_0_0_7/syncx_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_7/n287_q_reg[4]  ( .D(\fadd_0_0_0_0_7/syncx_d1 [4]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_7/syncx_d2 [4]) );
  DFFX1 \p_val_203_reg[4]  ( .D(n12580), .CLK(clk), .Q(n14010) );
  DFFX1 \p_val_294_reg[4]  ( .D(n12579), .CLK(clk), .Q(n13858) );
  DFFX1 \fadd_0_0_0_0_6_y_reg[4]  ( .D(n13011), .CLK(clk), .Q(n5550), .QN(
        n14601) );
  DFFX1 \fadd_0_0_0_0_7_x_reg[4]  ( .D(n13023), .CLK(clk), .Q(n5490), .QN(
        n14617) );
  DFFX1 \fadd_0_0_0_0_7/n275_q_reg[5]  ( .D(\fadd_0_0_0_0_7/newx [5]), .CLK(
        clk), .Q(\fadd_0_0_0_0_7/newx_d1 [5]) );
  DFFX1 \fadd_0_0_0_0_7/n281_q_reg[1]  ( .D(\fadd_0_0_0_0_7/newx [5]), .CLK(
        clk), .Q(\fadd_0_0_0_0_7/exponentresultfar0_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_7/n282_q_reg[1]  ( .D(
        \fadd_0_0_0_0_7/exponentresultfar0_d1 [1]), .CLK(clk), .Q(
        \fadd_0_0_0_0_7/exponentresultfar0_d2 [1]) );
  DFFX1 \fadd_0_0_0_0_7/n286_q_reg[5]  ( .D(\fadd_0_0_0_0_7/newx [5]), .CLK(
        clk), .Q(\fadd_0_0_0_0_7/syncx_d1 [5]) );
  DFFX1 \fadd_0_0_0_0_7/n287_q_reg[5]  ( .D(\fadd_0_0_0_0_7/syncx_d1 [5]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_7/syncx_d2 [5]) );
  DFFX1 \p_val_203_reg[5]  ( .D(n12578), .CLK(clk), .Q(n14011) );
  DFFX1 \p_val_294_reg[5]  ( .D(n12577), .CLK(clk), .Q(n13881) );
  DFFX1 \fadd_0_0_0_0_6_y_reg[5]  ( .D(n13010), .CLK(clk), .Q(n5551), .QN(
        n14600) );
  DFFX1 \fadd_0_0_0_0_7_x_reg[5]  ( .D(n13022), .CLK(clk), .Q(n5491), .QN(
        n14616) );
  DFFX1 \fadd_0_0_0_0_7/n275_q_reg[6]  ( .D(\fadd_0_0_0_0_7/newx [6]), .CLK(
        clk), .Q(\fadd_0_0_0_0_7/newx_d1 [6]) );
  DFFX1 \fadd_0_0_0_0_7/n281_q_reg[2]  ( .D(\fadd_0_0_0_0_7/newx [6]), .CLK(
        clk), .Q(\fadd_0_0_0_0_7/exponentresultfar0_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_7/n282_q_reg[2]  ( .D(
        \fadd_0_0_0_0_7/exponentresultfar0_d1 [2]), .CLK(clk), .Q(
        \fadd_0_0_0_0_7/exponentresultfar0_d2 [2]) );
  DFFX1 \fadd_0_0_0_0_7/n286_q_reg[6]  ( .D(\fadd_0_0_0_0_7/newx [6]), .CLK(
        clk), .Q(\fadd_0_0_0_0_7/syncx_d1 [6]) );
  DFFX1 \fadd_0_0_0_0_7/n287_q_reg[6]  ( .D(\fadd_0_0_0_0_7/syncx_d1 [6]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_7/syncx_d2 [6]) );
  DFFX1 \p_val_203_reg[6]  ( .D(n12576), .CLK(clk), .Q(n14012) );
  DFFX1 \p_val_294_reg[6]  ( .D(n12575), .CLK(clk), .Q(n13856) );
  DFFX1 \fadd_0_0_0_0_6_y_reg[6]  ( .D(n13009), .CLK(clk), .Q(n5552), .QN(
        n14599) );
  DFFX1 \fadd_0_0_0_0_7_x_reg[6]  ( .D(n13021), .CLK(clk), .Q(n5492), .QN(
        n14615) );
  DFFX1 \fadd_0_0_0_0_7/n275_q_reg[7]  ( .D(\fadd_0_0_0_0_7/newx [7]), .CLK(
        clk), .Q(\fadd_0_0_0_0_7/newx_d1 [7]) );
  DFFX1 \fadd_0_0_0_0_7/n281_q_reg[3]  ( .D(\fadd_0_0_0_0_7/newx [7]), .CLK(
        clk), .Q(\fadd_0_0_0_0_7/exponentresultfar0_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_7/n282_q_reg[3]  ( .D(
        \fadd_0_0_0_0_7/exponentresultfar0_d1 [3]), .CLK(clk), .Q(
        \fadd_0_0_0_0_7/exponentresultfar0_d2 [3]) );
  DFFX1 \fadd_0_0_0_0_7/n286_q_reg[7]  ( .D(\fadd_0_0_0_0_7/newx [7]), .CLK(
        clk), .Q(\fadd_0_0_0_0_7/syncx_d1 [7]) );
  DFFX1 \fadd_0_0_0_0_7/n287_q_reg[7]  ( .D(\fadd_0_0_0_0_7/syncx_d1 [7]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_7/syncx_d2 [7]) );
  DFFX1 \p_val_203_reg[7]  ( .D(n12574), .CLK(clk), .Q(n14013) );
  DFFX1 \p_val_294_reg[7]  ( .D(n12573), .CLK(clk), .Q(n13882) );
  DFFX1 \fadd_0_0_0_0_6_y_reg[7]  ( .D(n13008), .CLK(clk), .Q(n5553), .QN(
        n14598) );
  DFFX1 \fadd_0_0_0_0_7_x_reg[7]  ( .D(n13020), .CLK(clk), .Q(n5493), .QN(
        n14614) );
  DFFX1 \fadd_0_0_0_0_7/n275_q_reg[8]  ( .D(\fadd_0_0_0_0_7/newx [8]), .CLK(
        clk), .Q(\fadd_0_0_0_0_7/newx_d1 [8]) );
  DFFX1 \fadd_0_0_0_0_7/n280_q_reg[0]  ( .D(
        \fadd_0_0_0_0_7/exponentresultclose [0]), .CLK(clk), .Q(
        \fadd_0_0_0_0_7/exponentresultclose_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_7/n280_q_reg[1]  ( .D(
        \fadd_0_0_0_0_7/exponentresultclose [1]), .CLK(clk), .Q(
        \fadd_0_0_0_0_7/exponentresultclose_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_7/n280_q_reg[2]  ( .D(
        \fadd_0_0_0_0_7/exponentresultclose [2]), .CLK(clk), .Q(
        \fadd_0_0_0_0_7/exponentresultclose_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_7/n280_q_reg[3]  ( .D(
        \fadd_0_0_0_0_7/exponentresultclose [3]), .CLK(clk), .Q(
        \fadd_0_0_0_0_7/exponentresultclose_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_7/n280_q_reg[4]  ( .D(
        \fadd_0_0_0_0_7/exponentresultclose [4]), .CLK(clk), .Q(
        \fadd_0_0_0_0_7/exponentresultclose_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_7/n280_q_reg[6]  ( .D(n13659), .CLK(clk), .Q(
        \fadd_0_0_0_0_7/exponentresultclose_d1 [6]) );
  DFFX1 \fadd_0_0_0_0_7/n280_q_reg[5]  ( .D(n13659), .CLK(clk), .Q(
        \fadd_0_0_0_0_7/exponentresultclose_d1 [5]) );
  DFFX1 \fadd_0_0_0_0_7/n281_q_reg[4]  ( .D(\fadd_0_0_0_0_7/newx [8]), .CLK(
        clk), .Q(\fadd_0_0_0_0_7/exponentresultfar0_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_7/n282_q_reg[4]  ( .D(
        \fadd_0_0_0_0_7/exponentresultfar0_d1 [4]), .CLK(clk), .Q(
        \fadd_0_0_0_0_7/exponentresultfar0_d2 [4]) );
  DFFX1 \fadd_0_0_0_0_7/n286_q_reg[8]  ( .D(\fadd_0_0_0_0_7/newx [8]), .CLK(
        clk), .Q(\fadd_0_0_0_0_7/syncx_d1 [8]) );
  DFFX1 \fadd_0_0_0_0_7/n287_q_reg[8]  ( .D(\fadd_0_0_0_0_7/syncx_d1 [8]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_7/syncx_d2 [8]) );
  DFFX1 \p_val_203_reg[8]  ( .D(n12572), .CLK(clk), .Q(n14014) );
  DFFX1 \p_val_294_reg[8]  ( .D(n12571), .CLK(clk), .Q(n13883) );
  DFFX1 \fadd_0_0_0_0_6_y_reg[8]  ( .D(n13007), .CLK(clk), .Q(n5554), .QN(
        n14597) );
  DFFX1 \fadd_0_0_0_0_7_x_reg[8]  ( .D(n13019), .CLK(clk), .Q(n5494), .QN(
        n14613) );
  DFFX1 \fadd_0_0_0_0_7/rightshiftercomponent/n413_q_reg[2]  ( .D(n14821), 
        .CLK(clk), .Q(\fadd_0_0_0_0_7/rightshiftercomponent/ps_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_7/rightshiftercomponent/n416_q_reg[1]  ( .D(
        \fadd_0_0_0_0_7/rightshiftercomponent/level2[1] ), .CLK(clk), .QN(
        n11578) );
  DFFX1 \fadd_0_0_0_0_7/rightshiftercomponent/n416_q_reg[0]  ( .D(n12761), 
        .CLK(clk), .QN(n11579) );
  DFFX1 \fadd_0_0_0_0_7/rightshiftercomponent/n413_q_reg[1]  ( .D(n14824), 
        .CLK(clk), .Q(\fadd_0_0_0_0_7/rightshiftercomponent/ps_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_7/rightshiftercomponent/n417_q_reg  ( .D(
        \fadd_0_0_0_0_7/rightshiftercomponent/n389_o ), .CLK(clk), .Q(n14951)
         );
  DFFX1 \fadd_0_0_0_0_7/rightshiftercomponent/n418_q_reg[0]  ( .D(n12760), 
        .CLK(clk), .Q(\fadd_0_0_0_0_7/rightshiftercomponent/level1_d1[0] ) );
  DFFX1 \fadd_0_0_0_0_7/rightshiftercomponent/n419_q_reg[0]  ( .D(
        \fadd_0_0_0_0_7/rightshiftercomponent/level1_d1[0] ), .CLK(clk), .Q(
        \fadd_0_0_0_0_7/rightshiftercomponent/level1_d2[0] ) );
  DFFX1 \fadd_0_0_0_0_7/rightshiftercomponent/n413_q_reg[0]  ( .D(n12759), 
        .CLK(clk), .Q(\fadd_0_0_0_0_7/rightshiftercomponent/ps_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_7/rightshiftercomponent/n414_q_reg[0]  ( .D(
        \fadd_0_0_0_0_7/rightshiftercomponent/ps_d1 [0]), .CLK(clk), .Q(
        \fadd_0_0_0_0_7/rightshiftercomponent/ps_d2[0] ) );
  DFFX1 \fadd_0_0_0_0_7/n293_q_reg[1]  ( .D(\fadd_0_0_0_0_7/newy_11 ), .CLK(
        clk), .Q(\fadd_0_0_0_0_7/syncexnxy_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_7/n294_q_reg[1]  ( .D(\fadd_0_0_0_0_7/syncexnxy_d1 [1]), 
        .CLK(clk), .QN(n12238) );
  DFFX1 \fadd_0_0_0_0_7/n278_q_reg  ( .D(n14820), .CLK(clk), .Q(
        \fadd_0_0_0_0_7/selectclosepath_d1 ), .QN(n11581) );
  DFFX1 \fadd_0_0_0_0_7/n283_q_reg  ( .D(\fadd_0_0_0_0_7/zerofromclose ), 
        .CLK(clk), .Q(\fadd_0_0_0_0_7/zerofromclose_d1 ) );
  DFFX1 \fadd_0_0_0_0_7/n290_q_reg  ( .D(\fadd_0_0_0_0_7/ressign ), .CLK(clk), 
        .Q(\fadd_0_0_0_0_7/syncressign_d1 ) );
  DFFX1 \fadd_0_0_0_0_7/n291_q_reg  ( .D(\fadd_0_0_0_0_7/syncressign_d1 ), 
        .CLK(clk), .QN(n12212) );
  DFFX1 \p_val_203_reg[9]  ( .D(n12570), .CLK(clk), .Q(n14015) );
  DFFX1 \p_val_294_reg[9]  ( .D(n12569), .CLK(clk), .Q(n14106), .QN(n12211) );
  DFFX1 \fadd_0_0_0_0_6_y_reg[9]  ( .D(n13006), .CLK(clk), .QN(n11770) );
  DFFX1 \fadd_0_0_0_0_6/n288_q_reg  ( .D(\fadd_0_0_0_0_6/newy_9 ), .CLK(clk), 
        .Q(\fadd_0_0_0_0_6/syncsigny_d1 ) );
  DFFX1 \fadd_0_0_0_0_6/n289_q_reg  ( .D(\fadd_0_0_0_0_6/syncsigny_d1 ), .CLK(
        clk), .Q(\fadd_0_0_0_0_6/syncsigny_d2 ) );
  DFFX1 \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[7]  ( .D(
        n12754), .CLK(clk), .Q(
        \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [7]) );
  DFFX1 \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[7]  ( .D(
        \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [7]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [7]) );
  DFFX1 \fadd_0_0_0_0_6/n284_q_reg  ( .D(n12754), .CLK(clk), .Q(
        \fadd_0_0_0_0_6/synceffsub_d1 ) );
  DFFX1 \fadd_0_0_0_0_6/n285_q_reg  ( .D(\fadd_0_0_0_0_6/synceffsub_d1 ), 
        .CLK(clk), .QN(n12203) );
  DFFX1 \fadd_0_0_0_0_6/n276_q_reg  ( .D(n12754), .CLK(clk), .Q(
        \fadd_0_0_0_0_6/effsub_d1 ) );
  DFFX1 \fadd_0_0_0_0_6/n277_q_reg  ( .D(\fadd_0_0_0_0_6/effsub_d1 ), .CLK(clk), .QN(n11557) );
  DFFX1 \p_val_179_reg[11]  ( .D(n12568), .CLK(clk), .Q(n13929) );
  DFFX1 \p_val_293_reg[11]  ( .D(n12567), .CLK(clk), .Q(n13859) );
  DFFX1 \fadd_0_0_0_0_6_x_reg[11]  ( .D(n12992), .CLK(clk), .Q(n13508), .QN(
        n12757) );
  DFFX1 \fadd_0_0_0_0_6/n293_q_reg[3]  ( .D(\fadd_0_0_0_0_6/newx [11]), .CLK(
        clk), .Q(\fadd_0_0_0_0_6/syncexnxy_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_6/n294_q_reg[3]  ( .D(\fadd_0_0_0_0_6/syncexnxy_d1 [3]), 
        .CLK(clk), .Q(n13777), .QN(n12209) );
  DFFX1 \fadd_0_0_0_0_4_y_reg[11]  ( .D(n12980), .CLK(clk), .Q(n13621), .QN(
        n12736) );
  DFFX1 \p_val_179_reg[10]  ( .D(n12566), .CLK(clk), .Q(n13930) );
  DFFX1 \p_val_293_reg[10]  ( .D(n12565), .CLK(clk), .Q(n13860) );
  DFFX1 \fadd_0_0_0_0_6_x_reg[10]  ( .D(n12993), .CLK(clk), .Q(n13473), .QN(
        n12758) );
  DFFX1 \fadd_0_0_0_0_6/n293_q_reg[2]  ( .D(\fadd_0_0_0_0_6/newx [10]), .CLK(
        clk), .Q(\fadd_0_0_0_0_6/syncexnxy_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_6/n294_q_reg[2]  ( .D(\fadd_0_0_0_0_6/syncexnxy_d1 [2]), 
        .CLK(clk), .Q(n13728) );
  DFFX1 \fadd_0_0_0_0_6/n293_q_reg[0]  ( .D(\fadd_0_0_0_0_6/newy_10 ), .CLK(
        clk), .Q(\fadd_0_0_0_0_6/syncexnxy_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_6/n294_q_reg[0]  ( .D(\fadd_0_0_0_0_6/syncexnxy_d1 [0]), 
        .CLK(clk), .Q(n12208), .QN(n13746) );
  DFFX1 \fadd_0_0_0_0_6/n293_q_reg[1]  ( .D(\fadd_0_0_0_0_6/newy_11 ), .CLK(
        clk), .Q(\fadd_0_0_0_0_6/syncexnxy_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_6/n294_q_reg[1]  ( .D(\fadd_0_0_0_0_6/syncexnxy_d1 [1]), 
        .CLK(clk), .QN(n12207) );
  DFFX1 \p_val_179_reg[3]  ( .D(n12564), .CLK(clk), .Q(n13931) );
  DFFX1 \p_val_293_reg[3]  ( .D(n12563), .CLK(clk), .Q(n13861) );
  DFFX1 \fadd_0_0_0_0_6_x_reg[3]  ( .D(n13000), .CLK(clk), .Q(n13496), .QN(
        n11775) );
  DFFX1 \fadd_0_0_0_0_6/n286_q_reg[3]  ( .D(
        \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ), .CLK(clk), .Q(\fadd_0_0_0_0_6/syncx_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_6/n287_q_reg[3]  ( .D(\fadd_0_0_0_0_6/syncx_d1 [3]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_6/syncx_d2 [3]) );
  DFFX1 \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/n432_q_reg[5]  ( .D(
        \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ), .CLK(clk), .Q(\fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [5]) );
  DFFX1 \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/n433_q_reg[5]  ( .D(
        \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [5]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/x_d2 [5]) );
  DFFX1 \fadd_0_0_0_0_4_y_reg[3]  ( .D(n12988), .CLK(clk), .Q(n13707), .QN(
        n11785) );
  DFFX1 \p_val_179_reg[4]  ( .D(n12562), .CLK(clk), .Q(n13932) );
  DFFX1 \p_val_293_reg[4]  ( .D(n12561), .CLK(clk), .Q(n13862) );
  DFFX1 \fadd_0_0_0_0_6_x_reg[4]  ( .D(n12999), .CLK(clk), .Q(n5562), .QN(
        n14606) );
  DFFX1 \fadd_0_0_0_0_6/n275_q_reg[4]  ( .D(\fadd_0_0_0_0_6/newx [4]), .CLK(
        clk), .Q(\fadd_0_0_0_0_6/newx_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_6/n281_q_reg[0]  ( .D(\fadd_0_0_0_0_6/newx [4]), .CLK(
        clk), .Q(\fadd_0_0_0_0_6/exponentresultfar0_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_6/n282_q_reg[0]  ( .D(
        \fadd_0_0_0_0_6/exponentresultfar0_d1 [0]), .CLK(clk), .Q(
        \fadd_0_0_0_0_6/exponentresultfar0_d2 [0]) );
  DFFX1 \fadd_0_0_0_0_6/n286_q_reg[4]  ( .D(\fadd_0_0_0_0_6/newx [4]), .CLK(
        clk), .Q(\fadd_0_0_0_0_6/syncx_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_6/n287_q_reg[4]  ( .D(\fadd_0_0_0_0_6/syncx_d1 [4]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_6/syncx_d2 [4]) );
  DFFX1 \fadd_0_0_0_0_4_y_reg[4]  ( .D(n12987), .CLK(clk), .Q(n5694), .QN(
        n14579) );
  DFFX1 \p_val_179_reg[5]  ( .D(n12560), .CLK(clk), .Q(n13933) );
  DFFX1 \p_val_293_reg[5]  ( .D(n12559), .CLK(clk), .Q(n13863) );
  DFFX1 \fadd_0_0_0_0_6_x_reg[5]  ( .D(n12998), .CLK(clk), .Q(n5563), .QN(
        n14605) );
  DFFX1 \fadd_0_0_0_0_6/n275_q_reg[5]  ( .D(\fadd_0_0_0_0_6/newx [5]), .CLK(
        clk), .Q(\fadd_0_0_0_0_6/newx_d1 [5]) );
  DFFX1 \fadd_0_0_0_0_6/n281_q_reg[1]  ( .D(\fadd_0_0_0_0_6/newx [5]), .CLK(
        clk), .Q(\fadd_0_0_0_0_6/exponentresultfar0_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_6/n282_q_reg[1]  ( .D(
        \fadd_0_0_0_0_6/exponentresultfar0_d1 [1]), .CLK(clk), .Q(
        \fadd_0_0_0_0_6/exponentresultfar0_d2 [1]) );
  DFFX1 \fadd_0_0_0_0_6/n286_q_reg[5]  ( .D(\fadd_0_0_0_0_6/newx [5]), .CLK(
        clk), .Q(\fadd_0_0_0_0_6/syncx_d1 [5]) );
  DFFX1 \fadd_0_0_0_0_6/n287_q_reg[5]  ( .D(\fadd_0_0_0_0_6/syncx_d1 [5]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_6/syncx_d2 [5]) );
  DFFX1 \fadd_0_0_0_0_4_y_reg[5]  ( .D(n12986), .CLK(clk), .Q(n5695), .QN(
        n14578) );
  DFFX1 \p_val_179_reg[6]  ( .D(n12558), .CLK(clk), .Q(n13934) );
  DFFX1 \p_val_293_reg[6]  ( .D(n12557), .CLK(clk), .Q(n13864) );
  DFFX1 \fadd_0_0_0_0_6_x_reg[6]  ( .D(n12997), .CLK(clk), .Q(n5564), .QN(
        n14604) );
  DFFX1 \fadd_0_0_0_0_6/n275_q_reg[6]  ( .D(\fadd_0_0_0_0_6/newx [6]), .CLK(
        clk), .Q(\fadd_0_0_0_0_6/newx_d1 [6]) );
  DFFX1 \fadd_0_0_0_0_6/n281_q_reg[2]  ( .D(\fadd_0_0_0_0_6/newx [6]), .CLK(
        clk), .Q(\fadd_0_0_0_0_6/exponentresultfar0_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_6/n282_q_reg[2]  ( .D(
        \fadd_0_0_0_0_6/exponentresultfar0_d1 [2]), .CLK(clk), .Q(
        \fadd_0_0_0_0_6/exponentresultfar0_d2 [2]) );
  DFFX1 \fadd_0_0_0_0_6/n286_q_reg[6]  ( .D(\fadd_0_0_0_0_6/newx [6]), .CLK(
        clk), .Q(\fadd_0_0_0_0_6/syncx_d1 [6]) );
  DFFX1 \fadd_0_0_0_0_6/n287_q_reg[6]  ( .D(\fadd_0_0_0_0_6/syncx_d1 [6]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_6/syncx_d2 [6]) );
  DFFX1 \fadd_0_0_0_0_4_y_reg[6]  ( .D(n12985), .CLK(clk), .Q(n5696), .QN(
        n14577) );
  DFFX1 \p_val_179_reg[7]  ( .D(n12556), .CLK(clk), .Q(n13935) );
  DFFX1 \p_val_293_reg[7]  ( .D(n12555), .CLK(clk), .Q(n13865) );
  DFFX1 \fadd_0_0_0_0_6_x_reg[7]  ( .D(n12996), .CLK(clk), .Q(n5565), .QN(
        n14603) );
  DFFX1 \fadd_0_0_0_0_6/n275_q_reg[7]  ( .D(\fadd_0_0_0_0_6/newx [7]), .CLK(
        clk), .Q(\fadd_0_0_0_0_6/newx_d1 [7]) );
  DFFX1 \fadd_0_0_0_0_6/n281_q_reg[3]  ( .D(\fadd_0_0_0_0_6/newx [7]), .CLK(
        clk), .Q(\fadd_0_0_0_0_6/exponentresultfar0_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_6/n282_q_reg[3]  ( .D(
        \fadd_0_0_0_0_6/exponentresultfar0_d1 [3]), .CLK(clk), .Q(
        \fadd_0_0_0_0_6/exponentresultfar0_d2 [3]) );
  DFFX1 \fadd_0_0_0_0_6/n286_q_reg[7]  ( .D(\fadd_0_0_0_0_6/newx [7]), .CLK(
        clk), .Q(\fadd_0_0_0_0_6/syncx_d1 [7]) );
  DFFX1 \fadd_0_0_0_0_6/n287_q_reg[7]  ( .D(\fadd_0_0_0_0_6/syncx_d1 [7]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_6/syncx_d2 [7]) );
  DFFX1 \fadd_0_0_0_0_4_y_reg[7]  ( .D(n12984), .CLK(clk), .Q(n5697), .QN(
        n14576) );
  DFFX1 \p_val_179_reg[8]  ( .D(n12554), .CLK(clk), .Q(n13936) );
  DFFX1 \p_val_293_reg[8]  ( .D(n12553), .CLK(clk), .Q(n13866) );
  DFFX1 \fadd_0_0_0_0_6_x_reg[8]  ( .D(n12995), .CLK(clk), .Q(n5566), .QN(
        n14602) );
  DFFX1 \fadd_0_0_0_0_6/rightshiftercomponent/n413_q_reg[2]  ( .D(n14800), 
        .CLK(clk), .Q(\fadd_0_0_0_0_6/rightshiftercomponent/ps_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_6/rightshiftercomponent/n416_q_reg[1]  ( .D(
        \fadd_0_0_0_0_6/rightshiftercomponent/level2[1] ), .CLK(clk), .QN(
        n11565) );
  DFFX1 \fadd_0_0_0_0_6/rightshiftercomponent/n413_q_reg[1]  ( .D(n14803), 
        .CLK(clk), .Q(\fadd_0_0_0_0_6/rightshiftercomponent/ps_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[5]  ( .D(
        \fadd_0_0_0_0_6/fracyfarxorop [5]), .CLK(clk), .Q(
        \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [5]) );
  DFFX1 \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[5]  ( .D(
        \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [5]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [5]) );
  DFFX1 \fadd_0_0_0_0_6/rightshiftercomponent/n413_q_reg[0]  ( .D(n12751), 
        .CLK(clk), .Q(\fadd_0_0_0_0_6/rightshiftercomponent/ps_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_6/rightshiftercomponent/n414_q_reg[0]  ( .D(
        \fadd_0_0_0_0_6/rightshiftercomponent/ps_d1 [0]), .CLK(clk), .Q(
        \fadd_0_0_0_0_6/rightshiftercomponent/ps_d2[0] ) );
  DFFX1 \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[6]  ( .D(
        \fadd_0_0_0_0_6/fracyfarxorop [6]), .CLK(clk), .Q(
        \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [6]) );
  DFFX1 \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[6]  ( .D(
        \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [6]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [6]) );
  DFFX1 \fadd_0_0_0_0_6/n275_q_reg[8]  ( .D(\fadd_0_0_0_0_6/newx [8]), .CLK(
        clk), .Q(\fadd_0_0_0_0_6/newx_d1 [8]) );
  DFFX1 \fadd_0_0_0_0_6/n280_q_reg[0]  ( .D(
        \fadd_0_0_0_0_6/exponentresultclose [0]), .CLK(clk), .Q(
        \fadd_0_0_0_0_6/exponentresultclose_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_6/n280_q_reg[1]  ( .D(
        \fadd_0_0_0_0_6/exponentresultclose [1]), .CLK(clk), .Q(
        \fadd_0_0_0_0_6/exponentresultclose_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_6/n280_q_reg[2]  ( .D(
        \fadd_0_0_0_0_6/exponentresultclose [2]), .CLK(clk), .Q(
        \fadd_0_0_0_0_6/exponentresultclose_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_6/n280_q_reg[3]  ( .D(
        \fadd_0_0_0_0_6/exponentresultclose [3]), .CLK(clk), .Q(
        \fadd_0_0_0_0_6/exponentresultclose_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_6/n280_q_reg[4]  ( .D(
        \fadd_0_0_0_0_6/exponentresultclose [4]), .CLK(clk), .Q(
        \fadd_0_0_0_0_6/exponentresultclose_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_6/n280_q_reg[6]  ( .D(n13658), .CLK(clk), .Q(
        \fadd_0_0_0_0_6/exponentresultclose_d1 [6]) );
  DFFX1 \fadd_0_0_0_0_6/n280_q_reg[5]  ( .D(n13658), .CLK(clk), .Q(
        \fadd_0_0_0_0_6/exponentresultclose_d1 [5]) );
  DFFX1 \fadd_0_0_0_0_6/n281_q_reg[4]  ( .D(\fadd_0_0_0_0_6/newx [8]), .CLK(
        clk), .Q(\fadd_0_0_0_0_6/exponentresultfar0_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_6/n282_q_reg[4]  ( .D(
        \fadd_0_0_0_0_6/exponentresultfar0_d1 [4]), .CLK(clk), .Q(
        \fadd_0_0_0_0_6/exponentresultfar0_d2 [4]) );
  DFFX1 \fadd_0_0_0_0_6/n286_q_reg[8]  ( .D(\fadd_0_0_0_0_6/newx [8]), .CLK(
        clk), .Q(\fadd_0_0_0_0_6/syncx_d1 [8]) );
  DFFX1 \fadd_0_0_0_0_6/n287_q_reg[8]  ( .D(\fadd_0_0_0_0_6/syncx_d1 [8]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_6/syncx_d2 [8]) );
  DFFX1 \fadd_0_0_0_0_4_y_reg[8]  ( .D(n12983), .CLK(clk), .Q(n5698), .QN(
        n14575) );
  DFFX1 \p_val_179_reg[2]  ( .D(n12552), .CLK(clk), .Q(n13937) );
  DFFX1 \p_val_293_reg[2]  ( .D(n12551), .CLK(clk), .Q(n13867) );
  DFFX1 \fadd_0_0_0_0_6_x_reg[2]  ( .D(n13001), .CLK(clk), .Q(n13494), .QN(
        n11774) );
  DFFX1 \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[4]  ( .D(
        \fadd_0_0_0_0_6/fracyfarxorop [4]), .CLK(clk), .Q(
        \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[4]  ( .D(
        \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [4]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [4]) );
  DFFX1 \fadd_0_0_0_0_6/rightshiftercomponent/n416_q_reg[0]  ( .D(n12753), 
        .CLK(clk), .QN(n11566) );
  DFFX1 \fadd_0_0_0_0_6/n286_q_reg[2]  ( .D(
        \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ), .CLK(clk), .Q(\fadd_0_0_0_0_6/syncx_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_6/n287_q_reg[2]  ( .D(\fadd_0_0_0_0_6/syncx_d1 [2]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_6/syncx_d2 [2]) );
  DFFX1 \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/n432_q_reg[4]  ( .D(
        \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ), .CLK(clk), .Q(\fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/n433_q_reg[4]  ( .D(
        \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [4]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/x_d2 [4]) );
  DFFX1 \fadd_0_0_0_0_4_y_reg[2]  ( .D(n12989), .CLK(clk), .Q(n13685), .QN(
        n11784) );
  DFFX1 \p_val_179_reg[1]  ( .D(n12550), .CLK(clk), .Q(n13938) );
  DFFX1 \p_val_293_reg[1]  ( .D(n12549), .CLK(clk), .Q(n13868) );
  DFFX1 \fadd_0_0_0_0_6_x_reg[1]  ( .D(n13002), .CLK(clk), .Q(n13481), .QN(
        n11773) );
  DFFX1 \fadd_0_0_0_0_6/rightshiftercomponent/n415_q_reg[3]  ( .D(n14809), 
        .CLK(clk), .QN(n11564) );
  DFFX1 \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[3]  ( .D(
        \fadd_0_0_0_0_6/fracyfarxorop [3]), .CLK(clk), .Q(
        \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[3]  ( .D(
        \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [3]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [3]) );
  DFFX1 \fadd_0_0_0_0_6/n286_q_reg[1]  ( .D(
        \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ), .CLK(clk), .Q(\fadd_0_0_0_0_6/syncx_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_6/n287_q_reg[1]  ( .D(\fadd_0_0_0_0_6/syncx_d1 [1]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_6/syncx_d2 [1]) );
  DFFX1 \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/n432_q_reg[3]  ( .D(
        \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ), .CLK(clk), .Q(\fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/n433_q_reg[3]  ( .D(
        \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [3]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/x_d2 [3]) );
  DFFX1 \fadd_0_0_0_0_4_y_reg[1]  ( .D(n12990), .CLK(clk), .Q(n13664), .QN(
        n11783) );
  DFFX1 \p_val_179_reg[0]  ( .D(n12548), .CLK(clk), .Q(n13939) );
  DFFX1 \p_val_293_reg[0]  ( .D(n12547), .CLK(clk), .Q(n13869) );
  DFFX1 \fadd_0_0_0_0_6_x_reg[0]  ( .D(n13003), .CLK(clk), .Q(n13479), .QN(
        n11772) );
  DFFX1 \fadd_0_0_0_0_6/rightshiftercomponent/n415_q_reg[2]  ( .D(n14810), 
        .CLK(clk), .QN(n11563) );
  DFFX1 \fadd_0_0_0_0_6/rightshiftercomponent/n417_q_reg  ( .D(
        \fadd_0_0_0_0_6/rightshiftercomponent/n389_o ), .CLK(clk), .Q(n14953)
         );
  DFFX1 \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[2]  ( .D(
        \fadd_0_0_0_0_6/fracyfarxorop [2]), .CLK(clk), .Q(
        \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[2]  ( .D(
        \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [2]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [2]) );
  DFFX1 \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[1]  ( .D(
        \fadd_0_0_0_0_6/fracyfarxorop [1]), .CLK(clk), .Q(
        \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[1]  ( .D(
        \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [1]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [1]) );
  DFFX1 \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[0]  ( .D(
        \fadd_0_0_0_0_6/fracyfarxorop [0]), .CLK(clk), .Q(
        \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[0]  ( .D(
        \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [0]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [0]) );
  DFFX1 \fadd_0_0_0_0_6/rightshiftercomponent/n418_q_reg[0]  ( .D(n12752), 
        .CLK(clk), .Q(\fadd_0_0_0_0_6/rightshiftercomponent/level1_d1[0] ) );
  DFFX1 \fadd_0_0_0_0_6/rightshiftercomponent/n419_q_reg[0]  ( .D(
        \fadd_0_0_0_0_6/rightshiftercomponent/level1_d1[0] ), .CLK(clk), .Q(
        \fadd_0_0_0_0_6/rightshiftercomponent/level1_d2[0] ) );
  DFFX1 \fadd_0_0_0_0_6/n286_q_reg[0]  ( .D(
        \add_0_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .CLK(clk), .Q(\fadd_0_0_0_0_6/syncx_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_6/n287_q_reg[0]  ( .D(\fadd_0_0_0_0_6/syncx_d1 [0]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_6/syncx_d2 [0]) );
  DFFX1 \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/n432_q_reg[2]  ( .D(
        \add_0_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .CLK(clk), .Q(\fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/n433_q_reg[2]  ( .D(
        \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [2]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/x_d2 [2]) );
  DFFX1 \fadd_0_0_0_0_4_y_reg[0]  ( .D(n12991), .CLK(clk), .Q(n13636), .QN(
        n11782) );
  DFFX1 \fadd_0_0_0_0_6/n278_q_reg  ( .D(n14799), .CLK(clk), .Q(
        \fadd_0_0_0_0_6/selectclosepath_d1 ), .QN(n11568) );
  DFFX1 \fadd_0_0_0_0_6/n283_q_reg  ( .D(\fadd_0_0_0_0_6/zerofromclose ), 
        .CLK(clk), .Q(\fadd_0_0_0_0_6/zerofromclose_d1 ) );
  DFFX1 \fadd_0_0_0_0_6/n290_q_reg  ( .D(\fadd_0_0_0_0_6/ressign ), .CLK(clk), 
        .Q(\fadd_0_0_0_0_6/syncressign_d1 ) );
  DFFX1 \fadd_0_0_0_0_6/n291_q_reg  ( .D(\fadd_0_0_0_0_6/syncressign_d1 ), 
        .CLK(clk), .QN(n12182) );
  DFFX1 \p_val_179_reg[9]  ( .D(n12546), .CLK(clk), .Q(n13940) );
  DFFX1 \p_val_293_reg[9]  ( .D(n12545), .CLK(clk), .Q(n14107), .QN(n12181) );
  DFFX1 \fadd_0_0_0_0_6_x_reg[9]  ( .D(n12994), .CLK(clk), .QN(n11781) );
  DFFX1 \fadd_0_0_0_0_6/n286_q_reg[9]  ( .D(n14806), .CLK(clk), .Q(
        \fadd_0_0_0_0_6/syncx_d1 [9]) );
  DFFX1 \fadd_0_0_0_0_6/n287_q_reg[9]  ( .D(\fadd_0_0_0_0_6/syncx_d1 [9]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_6/syncx_d2 [9]) );
  DFFX1 \fadd_0_0_0_0_4_y_reg[9]  ( .D(n12982), .CLK(clk), .Q(n13716), .QN(
        n11791) );
  DFFX1 \fadd_0_0_0_0_4_y_reg[10]  ( .D(n12981), .CLK(clk), .Q(n13888), .QN(
        n11792) );
  DFFX1 \fadd_0_0_0_0_4/n293_q_reg[0]  ( .D(\fadd_0_0_0_0_4/newy_10 ), .CLK(
        clk), .Q(\fadd_0_0_0_0_4/syncexnxy_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_4/n294_q_reg[0]  ( .D(\fadd_0_0_0_0_4/syncexnxy_d1 [0]), 
        .CLK(clk), .Q(n12178) );
  DFFX1 \p_val_131_reg[9]  ( .D(n12544), .CLK(clk), .Q(n13816) );
  DFFX1 \p_val_291_reg[9]  ( .D(n12543), .CLK(clk), .Q(n13941) );
  DFFX1 \fadd_0_0_0_0_4_x_reg[9]  ( .D(n12970), .CLK(clk), .Q(n13584), .QN(
        n11802) );
  DFFX1 \fadd_0_0_0_0_4/n288_q_reg  ( .D(\fadd_0_0_0_0_4/newy_9 ), .CLK(clk), 
        .Q(\fadd_0_0_0_0_4/syncsigny_d1 ) );
  DFFX1 \fadd_0_0_0_0_4/n289_q_reg  ( .D(\fadd_0_0_0_0_4/syncsigny_d1 ), .CLK(
        clk), .QN(n12175) );
  DFFX1 \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[7]  ( .D(
        n12734), .CLK(clk), .Q(
        \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [7]) );
  DFFX1 \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[7]  ( .D(
        \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [7]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [7]) );
  DFFX1 \fadd_0_0_0_0_4/n284_q_reg  ( .D(n12734), .CLK(clk), .Q(
        \fadd_0_0_0_0_4/synceffsub_d1 ) );
  DFFX1 \fadd_0_0_0_0_4/n285_q_reg  ( .D(\fadd_0_0_0_0_4/synceffsub_d1 ), 
        .CLK(clk), .QN(n12169) );
  DFFX1 \fadd_0_0_0_0_4/n276_q_reg  ( .D(n12734), .CLK(clk), .Q(
        \fadd_0_0_0_0_4/effsub_d1 ) );
  DFFX1 \fadd_0_0_0_0_4/n277_q_reg  ( .D(\fadd_0_0_0_0_4/effsub_d1 ), .CLK(clk), .QN(n11531) );
  DFFX1 \p_val_131_reg[11]  ( .D(n12542), .CLK(clk), .Q(n13817) );
  DFFX1 \p_val_291_reg[11]  ( .D(n12541), .CLK(clk), .Q(n13942) );
  DFFX1 \fadd_0_0_0_0_4_x_reg[11]  ( .D(n12968), .CLK(clk), .Q(n13514), .QN(
        n12737) );
  DFFX1 \fadd_0_0_0_0_4/n293_q_reg[3]  ( .D(\fadd_0_0_0_0_4/newx [11]), .CLK(
        clk), .Q(\fadd_0_0_0_0_4/syncexnxy_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_4/n294_q_reg[3]  ( .D(\fadd_0_0_0_0_4/syncexnxy_d1 [3]), 
        .CLK(clk), .QN(n12176) );
  DFFX1 \fadd_0_0_0_0_0_y_reg[11]  ( .D(n12956), .CLK(clk), .Q(n13627), .QN(
        n12696) );
  DFFX1 \p_val_131_reg[10]  ( .D(n12540), .CLK(clk), .Q(n13818) );
  DFFX1 \p_val_291_reg[10]  ( .D(n12539), .CLK(clk), .Q(n13943) );
  DFFX1 \fadd_0_0_0_0_4_x_reg[10]  ( .D(n12969), .CLK(clk), .Q(n13505), .QN(
        n12738) );
  DFFX1 \fadd_0_0_0_0_4/n286_q_reg[9]  ( .D(n14753), .CLK(clk), .Q(
        \fadd_0_0_0_0_4/syncx_d1 [9]) );
  DFFX1 \fadd_0_0_0_0_4/n287_q_reg[9]  ( .D(\fadd_0_0_0_0_4/syncx_d1 [9]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_4/syncx_d2 [9]) );
  DFFX1 \fadd_0_0_0_0_4/n286_q_reg[0]  ( .D(
        \add_0_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .CLK(clk), .Q(\fadd_0_0_0_0_4/syncx_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_4/n287_q_reg[0]  ( .D(\fadd_0_0_0_0_4/syncx_d1 [0]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_4/syncx_d2 [0]) );
  DFFX1 \p_val_131_reg[0]  ( .D(n12538), .CLK(clk), .Q(n13819) );
  DFFX1 \p_val_291_reg[0]  ( .D(n12537), .CLK(clk), .Q(n13944) );
  DFFX1 \fadd_0_0_0_0_4_x_reg[0]  ( .D(n12979), .CLK(clk), .Q(n13522), .QN(
        n11793) );
  DFFX1 \fadd_0_0_0_0_4/rightshiftercomponent/n415_q_reg[2]  ( .D(n14757), 
        .CLK(clk), .QN(n11537) );
  DFFX1 \fadd_0_0_0_0_0_y_reg[0]  ( .D(n12967), .CLK(clk), .Q(n13642), .QN(
        n11803) );
  DFFX1 \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/n432_q_reg[2]  ( .D(
        \add_0_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .CLK(clk), .Q(\fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/n433_q_reg[2]  ( .D(
        \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [2]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/x_d2 [2]) );
  DFFX1 \fadd_0_0_0_0_4/n293_q_reg[2]  ( .D(\fadd_0_0_0_0_4/newx [10]), .CLK(
        clk), .Q(\fadd_0_0_0_0_4/syncexnxy_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_4/n294_q_reg[2]  ( .D(\fadd_0_0_0_0_4/syncexnxy_d1 [2]), 
        .CLK(clk), .Q(n13725), .QN(n12174) );
  DFFX1 \fadd_0_0_0_0_4/n286_q_reg[1]  ( .D(
        \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ), .CLK(clk), .Q(\fadd_0_0_0_0_4/syncx_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_4/n287_q_reg[1]  ( .D(\fadd_0_0_0_0_4/syncx_d1 [1]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_4/syncx_d2 [1]) );
  DFFX1 \p_val_131_reg[1]  ( .D(n12536), .CLK(clk), .Q(n13820) );
  DFFX1 \p_val_291_reg[1]  ( .D(n12535), .CLK(clk), .Q(n13945) );
  DFFX1 \fadd_0_0_0_0_4_x_reg[1]  ( .D(n12978), .CLK(clk), .Q(n13533), .QN(
        n11794) );
  DFFX1 \fadd_0_0_0_0_4/rightshiftercomponent/n415_q_reg[3]  ( .D(n14756), 
        .CLK(clk), .QN(n11538) );
  DFFX1 \fadd_0_0_0_0_0_y_reg[1]  ( .D(n12966), .CLK(clk), .Q(n13670), .QN(
        n11804) );
  DFFX1 \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/n432_q_reg[3]  ( .D(
        \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ), .CLK(clk), .Q(\fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/n433_q_reg[3]  ( .D(
        \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [3]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/x_d2 [3]) );
  DFFX1 \fadd_0_0_0_0_4/n286_q_reg[2]  ( .D(
        \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ), .CLK(clk), .Q(\fadd_0_0_0_0_4/syncx_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_4/n287_q_reg[2]  ( .D(\fadd_0_0_0_0_4/syncx_d1 [2]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_4/syncx_d2 [2]) );
  DFFX1 \p_val_131_reg[2]  ( .D(n12534), .CLK(clk), .Q(n13821) );
  DFFX1 \p_val_291_reg[2]  ( .D(n12533), .CLK(clk), .Q(n13946) );
  DFFX1 \fadd_0_0_0_0_4_x_reg[2]  ( .D(n12977), .CLK(clk), .Q(n13558), .QN(
        n11795) );
  DFFX1 \fadd_0_0_0_0_0_y_reg[2]  ( .D(n12965), .CLK(clk), .Q(n13691), .QN(
        n11805) );
  DFFX1 \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/n432_q_reg[4]  ( .D(
        \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ), .CLK(clk), .Q(\fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/n433_q_reg[4]  ( .D(
        \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [4]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/x_d2 [4]) );
  DFFX1 \fadd_0_0_0_0_4/n286_q_reg[3]  ( .D(
        \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ), .CLK(clk), .Q(\fadd_0_0_0_0_4/syncx_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_4/n287_q_reg[3]  ( .D(\fadd_0_0_0_0_4/syncx_d1 [3]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_4/syncx_d2 [3]) );
  DFFX1 \p_val_131_reg[3]  ( .D(n12532), .CLK(clk), .Q(n13822) );
  DFFX1 \p_val_291_reg[3]  ( .D(n12531), .CLK(clk), .Q(n13947) );
  DFFX1 \fadd_0_0_0_0_4_x_reg[3]  ( .D(n12976), .CLK(clk), .Q(n13575), .QN(
        n11796) );
  DFFX1 \fadd_0_0_0_0_0_y_reg[3]  ( .D(n12964), .CLK(clk), .Q(n13713), .QN(
        n11806) );
  DFFX1 \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/n432_q_reg[5]  ( .D(
        \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ), .CLK(clk), .Q(\fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [5]) );
  DFFX1 \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/n433_q_reg[5]  ( .D(
        \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [5]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/x_d2 [5]) );
  DFFX1 \fadd_0_0_0_0_4/n275_q_reg[4]  ( .D(\fadd_0_0_0_0_4/newx [4]), .CLK(
        clk), .Q(\fadd_0_0_0_0_4/newx_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_4/n281_q_reg[0]  ( .D(\fadd_0_0_0_0_4/newx [4]), .CLK(
        clk), .Q(\fadd_0_0_0_0_4/exponentresultfar0_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_4/n282_q_reg[0]  ( .D(
        \fadd_0_0_0_0_4/exponentresultfar0_d1 [0]), .CLK(clk), .Q(
        \fadd_0_0_0_0_4/exponentresultfar0_d2 [0]) );
  DFFX1 \fadd_0_0_0_0_4/n286_q_reg[4]  ( .D(\fadd_0_0_0_0_4/newx [4]), .CLK(
        clk), .Q(\fadd_0_0_0_0_4/syncx_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_4/n287_q_reg[4]  ( .D(\fadd_0_0_0_0_4/syncx_d1 [4]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_4/syncx_d2 [4]) );
  DFFX1 \p_val_131_reg[4]  ( .D(n12530), .CLK(clk), .Q(n13823) );
  DFFX1 \p_val_291_reg[4]  ( .D(n12529), .CLK(clk), .Q(n13948) );
  DFFX1 \fadd_0_0_0_0_4_x_reg[4]  ( .D(n12975), .CLK(clk), .Q(n5706), .QN(
        n14584) );
  DFFX1 \fadd_0_0_0_0_0_y_reg[4]  ( .D(n12963), .CLK(clk), .Q(n5982), .QN(
        n14535) );
  DFFX1 \fadd_0_0_0_0_4/n275_q_reg[5]  ( .D(\fadd_0_0_0_0_4/newx [5]), .CLK(
        clk), .Q(\fadd_0_0_0_0_4/newx_d1 [5]) );
  DFFX1 \fadd_0_0_0_0_4/n281_q_reg[1]  ( .D(\fadd_0_0_0_0_4/newx [5]), .CLK(
        clk), .Q(\fadd_0_0_0_0_4/exponentresultfar0_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_4/n282_q_reg[1]  ( .D(
        \fadd_0_0_0_0_4/exponentresultfar0_d1 [1]), .CLK(clk), .Q(
        \fadd_0_0_0_0_4/exponentresultfar0_d2 [1]) );
  DFFX1 \fadd_0_0_0_0_4/n286_q_reg[5]  ( .D(\fadd_0_0_0_0_4/newx [5]), .CLK(
        clk), .Q(\fadd_0_0_0_0_4/syncx_d1 [5]) );
  DFFX1 \fadd_0_0_0_0_4/n287_q_reg[5]  ( .D(\fadd_0_0_0_0_4/syncx_d1 [5]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_4/syncx_d2 [5]) );
  DFFX1 \p_val_131_reg[5]  ( .D(n12528), .CLK(clk), .Q(n13824) );
  DFFX1 \p_val_291_reg[5]  ( .D(n12527), .CLK(clk), .Q(n13949) );
  DFFX1 \fadd_0_0_0_0_4_x_reg[5]  ( .D(n12974), .CLK(clk), .Q(n5707), .QN(
        n14583) );
  DFFX1 \fadd_0_0_0_0_0_y_reg[5]  ( .D(n12962), .CLK(clk), .Q(n5983), .QN(
        n14534) );
  DFFX1 \fadd_0_0_0_0_4/n275_q_reg[6]  ( .D(\fadd_0_0_0_0_4/newx [6]), .CLK(
        clk), .Q(\fadd_0_0_0_0_4/newx_d1 [6]) );
  DFFX1 \fadd_0_0_0_0_4/n281_q_reg[2]  ( .D(\fadd_0_0_0_0_4/newx [6]), .CLK(
        clk), .Q(\fadd_0_0_0_0_4/exponentresultfar0_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_4/n282_q_reg[2]  ( .D(
        \fadd_0_0_0_0_4/exponentresultfar0_d1 [2]), .CLK(clk), .Q(
        \fadd_0_0_0_0_4/exponentresultfar0_d2 [2]) );
  DFFX1 \fadd_0_0_0_0_4/n286_q_reg[6]  ( .D(\fadd_0_0_0_0_4/newx [6]), .CLK(
        clk), .Q(\fadd_0_0_0_0_4/syncx_d1 [6]) );
  DFFX1 \fadd_0_0_0_0_4/n287_q_reg[6]  ( .D(\fadd_0_0_0_0_4/syncx_d1 [6]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_4/syncx_d2 [6]) );
  DFFX1 \p_val_131_reg[6]  ( .D(n12526), .CLK(clk), .Q(n13825) );
  DFFX1 \p_val_291_reg[6]  ( .D(n12525), .CLK(clk), .Q(n13950) );
  DFFX1 \fadd_0_0_0_0_4_x_reg[6]  ( .D(n12973), .CLK(clk), .Q(n5708), .QN(
        n14582) );
  DFFX1 \fadd_0_0_0_0_0_y_reg[6]  ( .D(n12961), .CLK(clk), .Q(n5984), .QN(
        n14533) );
  DFFX1 \fadd_0_0_0_0_4/n275_q_reg[7]  ( .D(\fadd_0_0_0_0_4/newx [7]), .CLK(
        clk), .Q(\fadd_0_0_0_0_4/newx_d1 [7]) );
  DFFX1 \fadd_0_0_0_0_4/n281_q_reg[3]  ( .D(\fadd_0_0_0_0_4/newx [7]), .CLK(
        clk), .Q(\fadd_0_0_0_0_4/exponentresultfar0_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_4/n282_q_reg[3]  ( .D(
        \fadd_0_0_0_0_4/exponentresultfar0_d1 [3]), .CLK(clk), .Q(
        \fadd_0_0_0_0_4/exponentresultfar0_d2 [3]) );
  DFFX1 \fadd_0_0_0_0_4/n286_q_reg[7]  ( .D(\fadd_0_0_0_0_4/newx [7]), .CLK(
        clk), .Q(\fadd_0_0_0_0_4/syncx_d1 [7]) );
  DFFX1 \fadd_0_0_0_0_4/n287_q_reg[7]  ( .D(\fadd_0_0_0_0_4/syncx_d1 [7]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_4/syncx_d2 [7]) );
  DFFX1 \p_val_131_reg[7]  ( .D(n12524), .CLK(clk), .Q(n13826) );
  DFFX1 \p_val_291_reg[7]  ( .D(n12523), .CLK(clk), .Q(n13951) );
  DFFX1 \fadd_0_0_0_0_4_x_reg[7]  ( .D(n12972), .CLK(clk), .Q(n5709), .QN(
        n14581) );
  DFFX1 \fadd_0_0_0_0_0_y_reg[7]  ( .D(n12960), .CLK(clk), .Q(n5985), .QN(
        n14532) );
  DFFX1 \fadd_0_0_0_0_4/n275_q_reg[8]  ( .D(\fadd_0_0_0_0_4/newx [8]), .CLK(
        clk), .Q(\fadd_0_0_0_0_4/newx_d1 [8]) );
  DFFX1 \fadd_0_0_0_0_4/n280_q_reg[0]  ( .D(
        \fadd_0_0_0_0_4/exponentresultclose [0]), .CLK(clk), .Q(
        \fadd_0_0_0_0_4/exponentresultclose_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_4/n280_q_reg[1]  ( .D(
        \fadd_0_0_0_0_4/exponentresultclose [1]), .CLK(clk), .Q(
        \fadd_0_0_0_0_4/exponentresultclose_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_4/n280_q_reg[2]  ( .D(
        \fadd_0_0_0_0_4/exponentresultclose [2]), .CLK(clk), .Q(
        \fadd_0_0_0_0_4/exponentresultclose_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_4/n280_q_reg[3]  ( .D(
        \fadd_0_0_0_0_4/exponentresultclose [3]), .CLK(clk), .Q(
        \fadd_0_0_0_0_4/exponentresultclose_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_4/n280_q_reg[4]  ( .D(
        \fadd_0_0_0_0_4/exponentresultclose [4]), .CLK(clk), .Q(
        \fadd_0_0_0_0_4/exponentresultclose_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_4/n280_q_reg[6]  ( .D(n13657), .CLK(clk), .Q(
        \fadd_0_0_0_0_4/exponentresultclose_d1 [6]) );
  DFFX1 \fadd_0_0_0_0_4/n280_q_reg[5]  ( .D(n13657), .CLK(clk), .Q(
        \fadd_0_0_0_0_4/exponentresultclose_d1 [5]) );
  DFFX1 \fadd_0_0_0_0_4/n281_q_reg[4]  ( .D(\fadd_0_0_0_0_4/newx [8]), .CLK(
        clk), .Q(\fadd_0_0_0_0_4/exponentresultfar0_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_4/n282_q_reg[4]  ( .D(
        \fadd_0_0_0_0_4/exponentresultfar0_d1 [4]), .CLK(clk), .Q(
        \fadd_0_0_0_0_4/exponentresultfar0_d2 [4]) );
  DFFX1 \fadd_0_0_0_0_4/n286_q_reg[8]  ( .D(\fadd_0_0_0_0_4/newx [8]), .CLK(
        clk), .Q(\fadd_0_0_0_0_4/syncx_d1 [8]) );
  DFFX1 \fadd_0_0_0_0_4/n287_q_reg[8]  ( .D(\fadd_0_0_0_0_4/syncx_d1 [8]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_4/syncx_d2 [8]) );
  DFFX1 \p_val_131_reg[8]  ( .D(n12522), .CLK(clk), .Q(n13827) );
  DFFX1 \p_val_291_reg[8]  ( .D(n12521), .CLK(clk), .Q(n13952) );
  DFFX1 \fadd_0_0_0_0_4_x_reg[8]  ( .D(n12971), .CLK(clk), .Q(n5710), .QN(
        n14580) );
  DFFX1 \fadd_0_0_0_0_4/rightshiftercomponent/n413_q_reg[2]  ( .D(n14747), 
        .CLK(clk), .Q(\fadd_0_0_0_0_4/rightshiftercomponent/ps_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_4/rightshiftercomponent/n416_q_reg[1]  ( .D(
        \fadd_0_0_0_0_4/rightshiftercomponent/level2[1] ), .CLK(clk), .QN(
        n11539) );
  DFFX1 \fadd_0_0_0_0_4/rightshiftercomponent/n416_q_reg[0]  ( .D(n12733), 
        .CLK(clk), .QN(n11540) );
  DFFX1 \fadd_0_0_0_0_4/rightshiftercomponent/n413_q_reg[1]  ( .D(n14750), 
        .CLK(clk), .Q(\fadd_0_0_0_0_4/rightshiftercomponent/ps_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_4/rightshiftercomponent/n417_q_reg  ( .D(
        \fadd_0_0_0_0_4/rightshiftercomponent/n389_o ), .CLK(clk), .Q(n14956)
         );
  DFFX1 \fadd_0_0_0_0_4/rightshiftercomponent/n418_q_reg[0]  ( .D(n12732), 
        .CLK(clk), .Q(\fadd_0_0_0_0_4/rightshiftercomponent/level1_d1[0] ) );
  DFFX1 \fadd_0_0_0_0_4/rightshiftercomponent/n419_q_reg[0]  ( .D(
        \fadd_0_0_0_0_4/rightshiftercomponent/level1_d1[0] ), .CLK(clk), .Q(
        \fadd_0_0_0_0_4/rightshiftercomponent/level1_d2[0] ) );
  DFFX1 \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[5]  ( .D(
        \fadd_0_0_0_0_4/fracyfarxorop [5]), .CLK(clk), .Q(
        \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [5]) );
  DFFX1 \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[5]  ( .D(
        \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [5]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [5]) );
  DFFX1 \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[3]  ( .D(
        \fadd_0_0_0_0_4/fracyfarxorop [3]), .CLK(clk), .Q(
        \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[3]  ( .D(
        \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [3]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [3]) );
  DFFX1 \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[2]  ( .D(
        \fadd_0_0_0_0_4/fracyfarxorop [2]), .CLK(clk), .Q(
        \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[2]  ( .D(
        \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [2]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [2]) );
  DFFX1 \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[1]  ( .D(
        \fadd_0_0_0_0_4/fracyfarxorop [1]), .CLK(clk), .Q(
        \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[1]  ( .D(
        \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [1]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [1]) );
  DFFX1 \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[0]  ( .D(
        \fadd_0_0_0_0_4/fracyfarxorop [0]), .CLK(clk), .Q(
        \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[0]  ( .D(
        \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [0]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [0]) );
  DFFX1 \fadd_0_0_0_0_4/rightshiftercomponent/n413_q_reg[0]  ( .D(n12731), 
        .CLK(clk), .Q(\fadd_0_0_0_0_4/rightshiftercomponent/ps_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_4/rightshiftercomponent/n414_q_reg[0]  ( .D(
        \fadd_0_0_0_0_4/rightshiftercomponent/ps_d1 [0]), .CLK(clk), .Q(
        \fadd_0_0_0_0_4/rightshiftercomponent/ps_d2[0] ) );
  DFFX1 \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[4]  ( .D(
        \fadd_0_0_0_0_4/fracyfarxorop [4]), .CLK(clk), .Q(
        \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[4]  ( .D(
        \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [4]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [4]) );
  DFFX1 \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[6]  ( .D(
        \fadd_0_0_0_0_4/fracyfarxorop [6]), .CLK(clk), .Q(
        \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [6]) );
  DFFX1 \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[6]  ( .D(
        \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [6]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [6]) );
  DFFX1 \fadd_0_0_0_0_0_y_reg[8]  ( .D(n12959), .CLK(clk), .Q(n5986), .QN(
        n14531) );
  DFFX1 \fadd_0_0_0_0_4/n293_q_reg[1]  ( .D(\fadd_0_0_0_0_4/newy_11 ), .CLK(
        clk), .Q(\fadd_0_0_0_0_4/syncexnxy_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_4/n294_q_reg[1]  ( .D(\fadd_0_0_0_0_4/syncexnxy_d1 [1]), 
        .CLK(clk), .Q(n13737), .QN(n12177) );
  DFFX1 \fadd_0_0_0_0_4/n278_q_reg  ( .D(n14746), .CLK(clk), .Q(
        \fadd_0_0_0_0_4/selectclosepath_d1 ), .QN(n11542) );
  DFFX1 \fadd_0_0_0_0_4/n283_q_reg  ( .D(\fadd_0_0_0_0_4/zerofromclose ), 
        .CLK(clk), .Q(\fadd_0_0_0_0_4/zerofromclose_d1 ) );
  DFFX1 \fadd_0_0_0_0_4/n290_q_reg  ( .D(\fadd_0_0_0_0_4/ressign ), .CLK(clk), 
        .Q(\fadd_0_0_0_0_4/syncressign_d1 ) );
  DFFX1 \fadd_0_0_0_0_4/n291_q_reg  ( .D(\fadd_0_0_0_0_4/syncressign_d1 ), 
        .CLK(clk), .QN(n12179) );
  DFFX1 \fadd_0_0_0_0_0_y_reg[10]  ( .D(n12957), .CLK(clk), .Q(n13894), .QN(
        n11813) );
  DFFX1 \fadd_0_0_0_0_0_y_reg[9]  ( .D(n12958), .CLK(clk), .QN(n11812) );
  DFFX1 \fadd_0_0_0_0_0/n288_q_reg  ( .D(\fadd_0_0_0_0_0/newy_9 ), .CLK(clk), 
        .Q(\fadd_0_0_0_0_0/syncsigny_d1 ) );
  DFFX1 \fadd_0_0_0_0_0/n289_q_reg  ( .D(\fadd_0_0_0_0_0/syncsigny_d1 ), .CLK(
        clk), .Q(\fadd_0_0_0_0_0/syncsigny_d2 ) );
  DFFX1 \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[7]  ( .D(
        n12694), .CLK(clk), .Q(
        \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [7]) );
  DFFX1 \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[7]  ( .D(
        \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [7]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [7]) );
  DFFX1 \fadd_0_0_0_0_0/n284_q_reg  ( .D(n12694), .CLK(clk), .Q(
        \fadd_0_0_0_0_0/synceffsub_d1 ) );
  DFFX1 \fadd_0_0_0_0_0/n285_q_reg  ( .D(\fadd_0_0_0_0_0/synceffsub_d1 ), 
        .CLK(clk), .QN(n12140) );
  DFFX1 \fadd_0_0_0_0_0/n276_q_reg  ( .D(n12694), .CLK(clk), .Q(
        \fadd_0_0_0_0_0/effsub_d1 ) );
  DFFX1 \fadd_0_0_0_0_0/n277_q_reg  ( .D(\fadd_0_0_0_0_0/effsub_d1 ), .CLK(clk), .QN(n11470) );
  DFFX1 \p_val_35_reg[11]  ( .D(n12520), .CLK(clk), .Q(n13828) );
  DFFX1 \p_val_287_reg[11]  ( .D(n12519), .CLK(clk), .Q(n13953) );
  DFFX1 \p_val_311_reg[11]  ( .D(n12518), .CLK(clk), .Q(n14094), .QN(n12142)
         );
  DFFX1 \fadd_0_0_0_0_0_x_reg[11]  ( .D(n12944), .CLK(clk), .Q(n13515), .QN(
        n12697) );
  DFFX1 \fadd_0_0_0_0_0/n293_q_reg[3]  ( .D(\fadd_0_0_0_0_0/newx [11]), .CLK(
        clk), .Q(\fadd_0_0_0_0_0/syncexnxy_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_0/n294_q_reg[3]  ( .D(\fadd_0_0_0_0_0/syncexnxy_d1 [3]), 
        .CLK(clk), .Q(n13778), .QN(n12148) );
  DFFX1 \p_val_35_reg[10]  ( .D(n12517), .CLK(clk), .Q(n13829) );
  DFFX1 \p_val_287_reg[10]  ( .D(n12516), .CLK(clk), .Q(n13954) );
  DFFX1 \p_val_311_reg[10]  ( .D(n12515), .CLK(clk), .Q(n14095), .QN(n12138)
         );
  DFFX1 \fadd_0_0_0_0_0_x_reg[10]  ( .D(n12945), .CLK(clk), .Q(n13506), .QN(
        n12698) );
  DFFX1 \fadd_0_0_0_0_0/n293_q_reg[2]  ( .D(\fadd_0_0_0_0_0/newx [10]), .CLK(
        clk), .Q(\fadd_0_0_0_0_0/syncexnxy_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_0/n294_q_reg[2]  ( .D(\fadd_0_0_0_0_0/syncexnxy_d1 [2]), 
        .CLK(clk), .Q(n13729) );
  DFFX1 \fadd_0_0_0_0_0/n293_q_reg[0]  ( .D(\fadd_0_0_0_0_0/newy_10 ), .CLK(
        clk), .Q(\fadd_0_0_0_0_0/syncexnxy_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_0/n294_q_reg[0]  ( .D(\fadd_0_0_0_0_0/syncexnxy_d1 [0]), 
        .CLK(clk), .Q(n12147), .QN(n13742) );
  DFFX1 \fadd_0_0_0_0_0/n293_q_reg[1]  ( .D(\fadd_0_0_0_0_0/newy_11 ), .CLK(
        clk), .Q(\fadd_0_0_0_0_0/syncexnxy_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_0/n294_q_reg[1]  ( .D(\fadd_0_0_0_0_0/syncexnxy_d1 [1]), 
        .CLK(clk), .QN(n12146) );
  DFFX1 \p_val_35_reg[0]  ( .D(n12514), .CLK(clk), .Q(n13830) );
  DFFX1 \p_val_287_reg[0]  ( .D(n12513), .CLK(clk), .Q(n13955) );
  DFFX1 \p_val_311_reg[0]  ( .D(n12512), .CLK(clk), .Q(n14096), .QN(n12135) );
  DFFX1 \fadd_0_0_0_0_0_x_reg[0]  ( .D(n12955), .CLK(clk), .Q(n13523), .QN(
        n11814) );
  DFFX1 \fadd_0_0_0_0_0/rightshiftercomponent/n415_q_reg[2]  ( .D(n14662), 
        .CLK(clk), .QN(n11476) );
  DFFX1 \fadd_0_0_0_0_0/n286_q_reg[0]  ( .D(
        \add_0_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .CLK(clk), .Q(\fadd_0_0_0_0_0/syncx_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_0/n287_q_reg[0]  ( .D(\fadd_0_0_0_0_0/syncx_d1 [0]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_0/syncx_d2 [0]) );
  DFFX1 \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/n432_q_reg[2]  ( .D(
        \add_0_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .CLK(clk), .Q(\fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/n433_q_reg[2]  ( .D(
        \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [2]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/x_d2 [2]) );
  DFFX1 \p_val_35_reg[1]  ( .D(n12511), .CLK(clk), .Q(n13831) );
  DFFX1 \p_val_287_reg[1]  ( .D(n12510), .CLK(clk), .Q(n13956) );
  DFFX1 \p_val_311_reg[1]  ( .D(n12509), .CLK(clk), .Q(n14097), .QN(n12132) );
  DFFX1 \fadd_0_0_0_0_0_x_reg[1]  ( .D(n12954), .CLK(clk), .Q(n13534), .QN(
        n11815) );
  DFFX1 \fadd_0_0_0_0_0/rightshiftercomponent/n415_q_reg[3]  ( .D(n14661), 
        .CLK(clk), .QN(n11477) );
  DFFX1 \fadd_0_0_0_0_0/n286_q_reg[1]  ( .D(
        \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ), .CLK(clk), .Q(\fadd_0_0_0_0_0/syncx_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_0/n287_q_reg[1]  ( .D(\fadd_0_0_0_0_0/syncx_d1 [1]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_0/syncx_d2 [1]) );
  DFFX1 \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/n432_q_reg[3]  ( .D(
        \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ), .CLK(clk), .Q(\fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/n433_q_reg[3]  ( .D(
        \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [3]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/x_d2 [3]) );
  DFFX1 \p_val_35_reg[2]  ( .D(n12508), .CLK(clk), .Q(n13832) );
  DFFX1 \p_val_287_reg[2]  ( .D(n12507), .CLK(clk), .Q(n13957) );
  DFFX1 \p_val_311_reg[2]  ( .D(n12506), .CLK(clk), .Q(n14098), .QN(n12129) );
  DFFX1 \fadd_0_0_0_0_0_x_reg[2]  ( .D(n12953), .CLK(clk), .Q(n13559), .QN(
        n11816) );
  DFFX1 \fadd_0_0_0_0_0/n286_q_reg[2]  ( .D(
        \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ), .CLK(clk), .Q(\fadd_0_0_0_0_0/syncx_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_0/n287_q_reg[2]  ( .D(\fadd_0_0_0_0_0/syncx_d1 [2]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_0/syncx_d2 [2]) );
  DFFX1 \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/n432_q_reg[4]  ( .D(
        \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ), .CLK(clk), .Q(\fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/n433_q_reg[4]  ( .D(
        \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [4]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/x_d2 [4]) );
  DFFX1 \p_val_35_reg[3]  ( .D(n12505), .CLK(clk), .Q(n13833) );
  DFFX1 \p_val_287_reg[3]  ( .D(n12504), .CLK(clk), .Q(n13958) );
  DFFX1 \p_val_311_reg[3]  ( .D(n12503), .CLK(clk), .Q(n14099), .QN(n12126) );
  DFFX1 \fadd_0_0_0_0_0_x_reg[3]  ( .D(n12952), .CLK(clk), .Q(n13576), .QN(
        n11817) );
  DFFX1 \fadd_0_0_0_0_0/n286_q_reg[3]  ( .D(
        \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ), .CLK(clk), .Q(\fadd_0_0_0_0_0/syncx_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_0/n287_q_reg[3]  ( .D(\fadd_0_0_0_0_0/syncx_d1 [3]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_0/syncx_d2 [3]) );
  DFFX1 \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/n432_q_reg[5]  ( .D(
        \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ), .CLK(clk), .Q(\fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [5]) );
  DFFX1 \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/n433_q_reg[5]  ( .D(
        \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [5]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/x_d2 [5]) );
  DFFX1 \p_val_35_reg[4]  ( .D(n12502), .CLK(clk), .Q(n13834) );
  DFFX1 \p_val_287_reg[4]  ( .D(n12501), .CLK(clk), .Q(n13959) );
  DFFX1 \p_val_311_reg[4]  ( .D(n12500), .CLK(clk), .Q(n14100), .QN(n12123) );
  DFFX1 \fadd_0_0_0_0_0_x_reg[4]  ( .D(n12951), .CLK(clk), .Q(n5994), .QN(
        n14540) );
  DFFX1 \fadd_0_0_0_0_0/n275_q_reg[4]  ( .D(\fadd_0_0_0_0_0/newx [4]), .CLK(
        clk), .Q(\fadd_0_0_0_0_0/newx_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_0/n281_q_reg[0]  ( .D(\fadd_0_0_0_0_0/newx [4]), .CLK(
        clk), .Q(\fadd_0_0_0_0_0/exponentresultfar0_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_0/n282_q_reg[0]  ( .D(
        \fadd_0_0_0_0_0/exponentresultfar0_d1 [0]), .CLK(clk), .Q(
        \fadd_0_0_0_0_0/exponentresultfar0_d2 [0]) );
  DFFX1 \fadd_0_0_0_0_0/n286_q_reg[4]  ( .D(\fadd_0_0_0_0_0/newx [4]), .CLK(
        clk), .Q(\fadd_0_0_0_0_0/syncx_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_0/n287_q_reg[4]  ( .D(\fadd_0_0_0_0_0/syncx_d1 [4]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_0/syncx_d2 [4]) );
  DFFX1 \p_val_35_reg[5]  ( .D(n12499), .CLK(clk), .Q(n13835) );
  DFFX1 \p_val_287_reg[5]  ( .D(n12498), .CLK(clk), .Q(n13960) );
  DFFX1 \p_val_311_reg[5]  ( .D(n12497), .CLK(clk), .Q(n14101), .QN(n12120) );
  DFFX1 \fadd_0_0_0_0_0_x_reg[5]  ( .D(n12950), .CLK(clk), .Q(n5995), .QN(
        n14539) );
  DFFX1 \fadd_0_0_0_0_0/n275_q_reg[5]  ( .D(\fadd_0_0_0_0_0/newx [5]), .CLK(
        clk), .Q(\fadd_0_0_0_0_0/newx_d1 [5]) );
  DFFX1 \fadd_0_0_0_0_0/n281_q_reg[1]  ( .D(\fadd_0_0_0_0_0/newx [5]), .CLK(
        clk), .Q(\fadd_0_0_0_0_0/exponentresultfar0_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_0/n282_q_reg[1]  ( .D(
        \fadd_0_0_0_0_0/exponentresultfar0_d1 [1]), .CLK(clk), .Q(
        \fadd_0_0_0_0_0/exponentresultfar0_d2 [1]) );
  DFFX1 \fadd_0_0_0_0_0/n286_q_reg[5]  ( .D(\fadd_0_0_0_0_0/newx [5]), .CLK(
        clk), .Q(\fadd_0_0_0_0_0/syncx_d1 [5]) );
  DFFX1 \fadd_0_0_0_0_0/n287_q_reg[5]  ( .D(\fadd_0_0_0_0_0/syncx_d1 [5]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_0/syncx_d2 [5]) );
  DFFX1 \p_val_35_reg[6]  ( .D(n12496), .CLK(clk), .Q(n13836) );
  DFFX1 \p_val_287_reg[6]  ( .D(n12495), .CLK(clk), .Q(n13961) );
  DFFX1 \p_val_311_reg[6]  ( .D(n12494), .CLK(clk), .Q(n14080), .QN(n12117) );
  DFFX1 \fadd_0_0_0_0_0_x_reg[6]  ( .D(n12949), .CLK(clk), .Q(n5996), .QN(
        n14538) );
  DFFX1 \fadd_0_0_0_0_0/n275_q_reg[6]  ( .D(\fadd_0_0_0_0_0/newx [6]), .CLK(
        clk), .Q(\fadd_0_0_0_0_0/newx_d1 [6]) );
  DFFX1 \fadd_0_0_0_0_0/n281_q_reg[2]  ( .D(\fadd_0_0_0_0_0/newx [6]), .CLK(
        clk), .Q(\fadd_0_0_0_0_0/exponentresultfar0_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_0/n282_q_reg[2]  ( .D(
        \fadd_0_0_0_0_0/exponentresultfar0_d1 [2]), .CLK(clk), .Q(
        \fadd_0_0_0_0_0/exponentresultfar0_d2 [2]) );
  DFFX1 \fadd_0_0_0_0_0/n286_q_reg[6]  ( .D(\fadd_0_0_0_0_0/newx [6]), .CLK(
        clk), .Q(\fadd_0_0_0_0_0/syncx_d1 [6]) );
  DFFX1 \fadd_0_0_0_0_0/n287_q_reg[6]  ( .D(\fadd_0_0_0_0_0/syncx_d1 [6]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_0/syncx_d2 [6]) );
  DFFX1 \p_val_35_reg[7]  ( .D(n12493), .CLK(clk), .Q(n13837) );
  DFFX1 \p_val_287_reg[7]  ( .D(n12492), .CLK(clk), .Q(n13962) );
  DFFX1 \p_val_311_reg[7]  ( .D(n12491), .CLK(clk), .Q(n14102), .QN(n12114) );
  DFFX1 \fadd_0_0_0_0_0_x_reg[7]  ( .D(n12948), .CLK(clk), .Q(n5997), .QN(
        n14537) );
  DFFX1 \fadd_0_0_0_0_0/n275_q_reg[7]  ( .D(\fadd_0_0_0_0_0/newx [7]), .CLK(
        clk), .Q(\fadd_0_0_0_0_0/newx_d1 [7]) );
  DFFX1 \fadd_0_0_0_0_0/n281_q_reg[3]  ( .D(\fadd_0_0_0_0_0/newx [7]), .CLK(
        clk), .Q(\fadd_0_0_0_0_0/exponentresultfar0_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_0/n282_q_reg[3]  ( .D(
        \fadd_0_0_0_0_0/exponentresultfar0_d1 [3]), .CLK(clk), .Q(
        \fadd_0_0_0_0_0/exponentresultfar0_d2 [3]) );
  DFFX1 \fadd_0_0_0_0_0/n286_q_reg[7]  ( .D(\fadd_0_0_0_0_0/newx [7]), .CLK(
        clk), .Q(\fadd_0_0_0_0_0/syncx_d1 [7]) );
  DFFX1 \fadd_0_0_0_0_0/n287_q_reg[7]  ( .D(\fadd_0_0_0_0_0/syncx_d1 [7]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_0/syncx_d2 [7]) );
  DFFX1 \p_val_35_reg[8]  ( .D(n12490), .CLK(clk), .Q(n13838) );
  DFFX1 \p_val_287_reg[8]  ( .D(n12489), .CLK(clk), .Q(n13963) );
  DFFX1 \p_val_311_reg[8]  ( .D(n12488), .CLK(clk), .Q(n14103), .QN(n12111) );
  DFFX1 \fadd_0_0_0_0_0_x_reg[8]  ( .D(n12947), .CLK(clk), .Q(n5998), .QN(
        n14536) );
  DFFX1 \fadd_0_0_0_0_0/rightshiftercomponent/n413_q_reg[2]  ( .D(n14652), 
        .CLK(clk), .Q(\fadd_0_0_0_0_0/rightshiftercomponent/ps_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_0/rightshiftercomponent/n416_q_reg[1]  ( .D(
        \fadd_0_0_0_0_0/rightshiftercomponent/level2[1] ), .CLK(clk), .QN(
        n11478) );
  DFFX1 \fadd_0_0_0_0_0/rightshiftercomponent/n416_q_reg[0]  ( .D(n12693), 
        .CLK(clk), .QN(n11479) );
  DFFX1 \fadd_0_0_0_0_0/rightshiftercomponent/n413_q_reg[1]  ( .D(n14655), 
        .CLK(clk), .Q(\fadd_0_0_0_0_0/rightshiftercomponent/ps_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_0/rightshiftercomponent/n417_q_reg  ( .D(
        \fadd_0_0_0_0_0/rightshiftercomponent/n389_o ), .CLK(clk), .Q(n14958)
         );
  DFFX1 \fadd_0_0_0_0_0/rightshiftercomponent/n418_q_reg[0]  ( .D(n12692), 
        .CLK(clk), .Q(\fadd_0_0_0_0_0/rightshiftercomponent/level1_d1[0] ) );
  DFFX1 \fadd_0_0_0_0_0/rightshiftercomponent/n419_q_reg[0]  ( .D(
        \fadd_0_0_0_0_0/rightshiftercomponent/level1_d1[0] ), .CLK(clk), .Q(
        \fadd_0_0_0_0_0/rightshiftercomponent/level1_d2[0] ) );
  DFFX1 \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[5]  ( .D(
        \fadd_0_0_0_0_0/fracyfarxorop [5]), .CLK(clk), .Q(
        \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [5]) );
  DFFX1 \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[5]  ( .D(
        \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [5]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [5]) );
  DFFX1 \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[3]  ( .D(
        \fadd_0_0_0_0_0/fracyfarxorop [3]), .CLK(clk), .Q(
        \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[3]  ( .D(
        \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [3]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [3]) );
  DFFX1 \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[2]  ( .D(
        \fadd_0_0_0_0_0/fracyfarxorop [2]), .CLK(clk), .Q(
        \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[2]  ( .D(
        \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [2]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [2]) );
  DFFX1 \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[1]  ( .D(
        \fadd_0_0_0_0_0/fracyfarxorop [1]), .CLK(clk), .Q(
        \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[1]  ( .D(
        \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [1]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [1]) );
  DFFX1 \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[0]  ( .D(
        \fadd_0_0_0_0_0/fracyfarxorop [0]), .CLK(clk), .Q(
        \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[0]  ( .D(
        \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [0]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [0]) );
  DFFX1 \fadd_0_0_0_0_0/rightshiftercomponent/n413_q_reg[0]  ( .D(n12691), 
        .CLK(clk), .Q(\fadd_0_0_0_0_0/rightshiftercomponent/ps_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_0/rightshiftercomponent/n414_q_reg[0]  ( .D(
        \fadd_0_0_0_0_0/rightshiftercomponent/ps_d1 [0]), .CLK(clk), .Q(
        \fadd_0_0_0_0_0/rightshiftercomponent/ps_d2[0] ) );
  DFFX1 \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[4]  ( .D(
        \fadd_0_0_0_0_0/fracyfarxorop [4]), .CLK(clk), .Q(
        \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[4]  ( .D(
        \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [4]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [4]) );
  DFFX1 \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[6]  ( .D(
        \fadd_0_0_0_0_0/fracyfarxorop [6]), .CLK(clk), .Q(
        \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [6]) );
  DFFX1 \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[6]  ( .D(
        \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [6]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [6]) );
  DFFX1 \fadd_0_0_0_0_0/n275_q_reg[8]  ( .D(\fadd_0_0_0_0_0/newx [8]), .CLK(
        clk), .Q(\fadd_0_0_0_0_0/newx_d1 [8]) );
  DFFX1 \fadd_0_0_0_0_0/n280_q_reg[0]  ( .D(
        \fadd_0_0_0_0_0/exponentresultclose [0]), .CLK(clk), .Q(
        \fadd_0_0_0_0_0/exponentresultclose_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_0/n280_q_reg[1]  ( .D(
        \fadd_0_0_0_0_0/exponentresultclose [1]), .CLK(clk), .Q(
        \fadd_0_0_0_0_0/exponentresultclose_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_0/n280_q_reg[2]  ( .D(
        \fadd_0_0_0_0_0/exponentresultclose [2]), .CLK(clk), .Q(
        \fadd_0_0_0_0_0/exponentresultclose_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_0/n280_q_reg[3]  ( .D(
        \fadd_0_0_0_0_0/exponentresultclose [3]), .CLK(clk), .Q(
        \fadd_0_0_0_0_0/exponentresultclose_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_0/n280_q_reg[4]  ( .D(
        \fadd_0_0_0_0_0/exponentresultclose [4]), .CLK(clk), .Q(
        \fadd_0_0_0_0_0/exponentresultclose_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_0/n280_q_reg[6]  ( .D(n13656), .CLK(clk), .Q(
        \fadd_0_0_0_0_0/exponentresultclose_d1 [6]) );
  DFFX1 \fadd_0_0_0_0_0/n280_q_reg[5]  ( .D(n13656), .CLK(clk), .Q(
        \fadd_0_0_0_0_0/exponentresultclose_d1 [5]) );
  DFFX1 \fadd_0_0_0_0_0/n281_q_reg[4]  ( .D(\fadd_0_0_0_0_0/newx [8]), .CLK(
        clk), .Q(\fadd_0_0_0_0_0/exponentresultfar0_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_0/n282_q_reg[4]  ( .D(
        \fadd_0_0_0_0_0/exponentresultfar0_d1 [4]), .CLK(clk), .Q(
        \fadd_0_0_0_0_0/exponentresultfar0_d2 [4]) );
  DFFX1 \fadd_0_0_0_0_0/n286_q_reg[8]  ( .D(\fadd_0_0_0_0_0/newx [8]), .CLK(
        clk), .Q(\fadd_0_0_0_0_0/syncx_d1 [8]) );
  DFFX1 \fadd_0_0_0_0_0/n287_q_reg[8]  ( .D(\fadd_0_0_0_0_0/syncx_d1 [8]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_0/syncx_d2 [8]) );
  DFFX1 \fadd_0_0_0_0_0/n278_q_reg  ( .D(n14651), .CLK(clk), .Q(
        \fadd_0_0_0_0_0/selectclosepath_d1 ), .QN(n11481) );
  DFFX1 \fadd_0_0_0_0_0/n283_q_reg  ( .D(\fadd_0_0_0_0_0/zerofromclose ), 
        .CLK(clk), .Q(\fadd_0_0_0_0_0/zerofromclose_d1 ) );
  DFFX1 \fadd_0_0_0_0_0/n290_q_reg  ( .D(\fadd_0_0_0_0_0/ressign ), .CLK(clk), 
        .Q(\fadd_0_0_0_0_0/syncressign_d1 ) );
  DFFX1 \fadd_0_0_0_0_0/n291_q_reg  ( .D(\fadd_0_0_0_0_0/syncressign_d1 ), 
        .CLK(clk), .QN(n12109) );
  DFFX1 \p_val_35_reg[9]  ( .D(n12487), .CLK(clk), .Q(n13839) );
  DFFX1 \p_val_287_reg[9]  ( .D(n12486), .CLK(clk), .Q(n13964) );
  DFFX1 \p_val_311_reg[9]  ( .D(n12485), .CLK(clk), .Q(n14104), .QN(n12107) );
  DFFX1 \fadd_0_0_0_0_0_x_reg[9]  ( .D(n12946), .CLK(clk), .Q(n13595), .QN(
        n11823) );
  DFFX1 \fadd_0_0_0_0_0/n286_q_reg[9]  ( .D(n14658), .CLK(clk), .Q(
        \fadd_0_0_0_0_0/syncx_d1 [9]) );
  DFFX1 \fadd_0_0_0_0_0/n287_q_reg[9]  ( .D(\fadd_0_0_0_0_0/syncx_d1 [9]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_0/syncx_d2 [9]) );
  DFFX1 \fadd_0_0_0_0_7_x_reg[9]  ( .D(n13018), .CLK(clk), .Q(n13582), .QN(
        n11760) );
  DFFX1 \fadd_0_0_0_0_7/n286_q_reg[9]  ( .D(n14827), .CLK(clk), .Q(
        \fadd_0_0_0_0_7/syncx_d1 [9]) );
  DFFX1 \fadd_0_0_0_0_7/n287_q_reg[9]  ( .D(\fadd_0_0_0_0_7/syncx_d1 [9]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_7/syncx_d2 [9]) );
  DFFX1 \fadd_0_0_0_0_7/n288_q_reg  ( .D(\fadd_0_0_0_0_7/newy_9 ), .CLK(clk), 
        .Q(\fadd_0_0_0_0_7/syncsigny_d1 ) );
  DFFX1 \fadd_0_0_0_0_7/n289_q_reg  ( .D(\fadd_0_0_0_0_7/syncsigny_d1 ), .CLK(
        clk), .Q(\fadd_0_0_0_0_7/syncsigny_d2 ) );
  DFFX1 \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[6]  ( .D(
        \fadd_0_0_0_0_7/fracyfarxorop [6]), .CLK(clk), .Q(
        \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [6]) );
  DFFX1 \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[6]  ( .D(
        \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [6]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [6]) );
  DFFX1 \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[4]  ( .D(
        \fadd_0_0_0_0_7/fracyfarxorop [4]), .CLK(clk), .Q(
        \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[4]  ( .D(
        \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [4]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [4]) );
  DFFX1 \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[3]  ( .D(
        \fadd_0_0_0_0_7/fracyfarxorop [3]), .CLK(clk), .Q(
        \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[3]  ( .D(
        \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [3]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [3]) );
  DFFX1 \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[2]  ( .D(
        \fadd_0_0_0_0_7/fracyfarxorop [2]), .CLK(clk), .Q(
        \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[2]  ( .D(
        \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [2]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [2]) );
  DFFX1 \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[1]  ( .D(
        \fadd_0_0_0_0_7/fracyfarxorop [1]), .CLK(clk), .Q(
        \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[1]  ( .D(
        \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [1]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [1]) );
  DFFX1 \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[0]  ( .D(
        \fadd_0_0_0_0_7/fracyfarxorop [0]), .CLK(clk), .Q(
        \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[0]  ( .D(
        \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [0]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [0]) );
  DFFX1 \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[5]  ( .D(
        \fadd_0_0_0_0_7/fracyfarxorop [5]), .CLK(clk), .Q(
        \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [5]) );
  DFFX1 \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[5]  ( .D(
        \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [5]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [5]) );
  DFFX1 \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[7]  ( .D(
        n12762), .CLK(clk), .Q(
        \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [7]) );
  DFFX1 \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[7]  ( .D(
        \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [7]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [7]) );
  DFFX1 \fadd_0_0_0_0_7/n284_q_reg  ( .D(n12762), .CLK(clk), .Q(
        \fadd_0_0_0_0_7/synceffsub_d1 ) );
  DFFX1 \fadd_0_0_0_0_7/n285_q_reg  ( .D(\fadd_0_0_0_0_7/synceffsub_d1 ), 
        .CLK(clk), .QN(n12231) );
  DFFX1 \fadd_0_0_0_0_7/n276_q_reg  ( .D(n12762), .CLK(clk), .Q(
        \fadd_0_0_0_0_7/effsub_d1 ) );
  DFFX1 \fadd_0_0_0_0_7/n277_q_reg  ( .D(\fadd_0_0_0_0_7/effsub_d1 ), .CLK(clk), .QN(n11570) );
  DFFX1 \fmul_0_0_0_0_8/roundingadder/n155_q_reg[0]  ( .D(
        \fmul_0_0_0_0_8/sigprodext [6]), .CLK(clk), .Q(
        \fmul_0_0_0_0_8/roundingadder/x_1_d1 [0]) );
  DFFX1 \fmul_0_0_0_0_8/roundingadder/n155_q_reg[1]  ( .D(
        \fmul_0_0_0_0_8/sigprodext [7]), .CLK(clk), .Q(
        \fmul_0_0_0_0_8/roundingadder/x_1_d1 [1]) );
  DFFX1 \fmul_0_0_0_0_8/roundingadder/n155_q_reg[2]  ( .D(
        \fmul_0_0_0_0_8/sigprodext [8]), .CLK(clk), .Q(
        \fmul_0_0_0_0_8/roundingadder/x_1_d1 [2]) );
  DFFX1 \fmul_0_0_0_0_8/roundingadder/n155_q_reg[3]  ( .D(
        \fmul_0_0_0_0_8/sigprodext [9]), .CLK(clk), .Q(
        \fmul_0_0_0_0_8/roundingadder/x_1_d1 [3]) );
  DFFX1 \fmul_0_0_0_0_8/roundingadder/n155_q_reg[4]  ( .D(
        \fmul_0_0_0_0_8/exppostnorm [0]), .CLK(clk), .Q(
        \fmul_0_0_0_0_8/roundingadder/x_1_d1 [4]) );
  DFFX1 \fmul_0_0_0_0_8/roundingadder/n155_q_reg[5]  ( .D(
        \fmul_0_0_0_0_8/exppostnorm [1]), .CLK(clk), .Q(
        \fmul_0_0_0_0_8/roundingadder/x_1_d1 [5]) );
  DFFX1 \fmul_0_0_0_0_8/roundingadder/n155_q_reg[6]  ( .D(
        \fmul_0_0_0_0_8/exppostnorm [2]), .CLK(clk), .Q(
        \fmul_0_0_0_0_8/roundingadder/x_1_d1 [6]) );
  DFFX1 \fmul_0_0_0_0_8/roundingadder/n155_q_reg[7]  ( .D(
        \fmul_0_0_0_0_8/exppostnorm [3]), .CLK(clk), .Q(
        \fmul_0_0_0_0_8/roundingadder/x_1_d1 [7]) );
  DFFX1 \fmul_0_0_0_0_8/roundingadder/n155_q_reg[8]  ( .D(
        \fmul_0_0_0_0_8/exppostnorm [4]), .CLK(clk), .Q(
        \fmul_0_0_0_0_8/roundingadder/x_1_d1 [8]) );
  DFFX1 \fmul_0_0_0_0_8/roundingadder/n155_q_reg[9]  ( .D(
        \fmul_0_0_0_0_8/exppostnorm [5]), .CLK(clk), .Q(
        \fmul_0_0_0_0_8/roundingadder/x_1_d1 [9]), .QN(n14170) );
  DFFX1 \fmul_0_0_0_0_8/roundingadder/n155_q_reg[10]  ( .D(n14129), .CLK(clk), 
        .Q(\fmul_0_0_0_0_8/roundingadder/x_1_d1 [10]) );
  DFFX1 \fmul_0_0_0_0_8/roundingadder/n154_q_reg  ( .D(\fmul_0_0_0_0_8/round ), 
        .CLK(clk), .Q(\fmul_0_0_0_0_8/roundingadder/n151_o[0] ) );
  DFFX1 \fmul_0_0_0_0_9/roundingadder/n155_q_reg[0]  ( .D(
        \fmul_0_0_0_0_9/sigprodext [6]), .CLK(clk), .Q(
        \fmul_0_0_0_0_9/roundingadder/x_1_d1 [0]) );
  DFFX1 \fmul_0_0_0_0_9/roundingadder/n155_q_reg[1]  ( .D(
        \fmul_0_0_0_0_9/sigprodext [7]), .CLK(clk), .Q(
        \fmul_0_0_0_0_9/roundingadder/x_1_d1 [1]) );
  DFFX1 \fmul_0_0_0_0_9/roundingadder/n155_q_reg[2]  ( .D(
        \fmul_0_0_0_0_9/sigprodext [8]), .CLK(clk), .Q(
        \fmul_0_0_0_0_9/roundingadder/x_1_d1 [2]) );
  DFFX1 \fmul_0_0_0_0_9/roundingadder/n155_q_reg[3]  ( .D(
        \fmul_0_0_0_0_9/sigprodext [9]), .CLK(clk), .Q(
        \fmul_0_0_0_0_9/roundingadder/x_1_d1 [3]) );
  DFFX1 \fmul_0_0_0_0_9/roundingadder/n155_q_reg[4]  ( .D(
        \fmul_0_0_0_0_9/exppostnorm [0]), .CLK(clk), .Q(
        \fmul_0_0_0_0_9/roundingadder/x_1_d1 [4]) );
  DFFX1 \fmul_0_0_0_0_9/roundingadder/n155_q_reg[5]  ( .D(
        \fmul_0_0_0_0_9/exppostnorm [1]), .CLK(clk), .Q(
        \fmul_0_0_0_0_9/roundingadder/x_1_d1 [5]) );
  DFFX1 \fmul_0_0_0_0_9/roundingadder/n155_q_reg[6]  ( .D(
        \fmul_0_0_0_0_9/exppostnorm [2]), .CLK(clk), .Q(
        \fmul_0_0_0_0_9/roundingadder/x_1_d1 [6]) );
  DFFX1 \fmul_0_0_0_0_9/roundingadder/n155_q_reg[7]  ( .D(
        \fmul_0_0_0_0_9/exppostnorm [3]), .CLK(clk), .Q(
        \fmul_0_0_0_0_9/roundingadder/x_1_d1 [7]) );
  DFFX1 \fmul_0_0_0_0_9/roundingadder/n155_q_reg[8]  ( .D(
        \fmul_0_0_0_0_9/exppostnorm [4]), .CLK(clk), .Q(
        \fmul_0_0_0_0_9/roundingadder/x_1_d1 [8]) );
  DFFX1 \fmul_0_0_0_0_9/roundingadder/n155_q_reg[9]  ( .D(
        \fmul_0_0_0_0_9/exppostnorm [5]), .CLK(clk), .Q(
        \fmul_0_0_0_0_9/roundingadder/x_1_d1 [9]) );
  DFFX1 \fmul_0_0_0_0_9/roundingadder/n155_q_reg[10]  ( .D(n14128), .CLK(clk), 
        .Q(\fmul_0_0_0_0_9/roundingadder/x_1_d1 [10]) );
  DFFX1 \fmul_0_0_0_0_9/roundingadder/n154_q_reg  ( .D(\fmul_0_0_0_0_9/round ), 
        .CLK(clk), .Q(\fmul_0_0_0_0_9/roundingadder/n151_o[0] ) );
  DFFX1 \fadd_0_0_0_0_9_y_reg[0]  ( .D(n12943), .CLK(clk), .Q(n13641), .QN(
        n11824) );
  DFFX1 \fadd_0_0_0_0_9_y_reg[1]  ( .D(n12942), .CLK(clk), .Q(n13669), .QN(
        n11825) );
  DFFX1 \fadd_0_0_0_0_9_y_reg[2]  ( .D(n12941), .CLK(clk), .Q(n13690), .QN(
        n11826) );
  DFFX1 \fadd_0_0_0_0_9_y_reg[3]  ( .D(n12940), .CLK(clk), .Q(n13712), .QN(
        n11827) );
  DFFX1 \fadd_0_0_0_0_9_y_reg[4]  ( .D(n12939), .CLK(clk), .Q(n5334), .QN(
        n14634) );
  DFFX1 \fadd_0_0_0_0_9_y_reg[5]  ( .D(n12938), .CLK(clk), .Q(n5335), .QN(
        n14633) );
  DFFX1 \fadd_0_0_0_0_9_y_reg[6]  ( .D(n12937), .CLK(clk), .Q(n5336), .QN(
        n14632) );
  DFFX1 \fadd_0_0_0_0_9_y_reg[7]  ( .D(n12936), .CLK(clk), .Q(n5337), .QN(
        n14631) );
  DFFX1 \fadd_0_0_0_0_9_y_reg[8]  ( .D(n12935), .CLK(clk), .Q(n5338), .QN(
        n14630) );
  DFFX1 \fadd_0_0_0_0_9_y_reg[11]  ( .D(n12932), .CLK(clk), .Q(n13626), .QN(
        n12786) );
  DFFX1 \fadd_0_0_0_0_9_y_reg[10]  ( .D(n12933), .CLK(clk), .Q(n13893), .QN(
        n11834) );
  DFFX1 \fadd_0_0_0_0_9/n293_q_reg[0]  ( .D(\fadd_0_0_0_0_9/newy_10 ), .CLK(
        clk), .Q(\fadd_0_0_0_0_9/syncexnxy_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_9/n294_q_reg[0]  ( .D(\fadd_0_0_0_0_9/syncexnxy_d1 [0]), 
        .CLK(clk), .Q(n12104) );
  DFFX1 \p_val_251_reg[9]  ( .D(n12484), .CLK(clk), .Q(n14016) );
  DFFX1 \p_val_296_reg[9]  ( .D(n12483), .CLK(clk), .Q(n14091), .QN(n12099) );
  DFFX1 \fadd_0_0_0_0_9_x_reg[9]  ( .D(n12922), .CLK(clk), .Q(n13583), .QN(
        n11844) );
  DFFX1 \fadd_0_0_0_0_9/n288_q_reg  ( .D(\fadd_0_0_0_0_9/newy_9 ), .CLK(clk), 
        .Q(\fadd_0_0_0_0_9/syncsigny_d1 ) );
  DFFX1 \fadd_0_0_0_0_9/n289_q_reg  ( .D(\fadd_0_0_0_0_9/syncsigny_d1 ), .CLK(
        clk), .QN(n12101) );
  DFFX1 \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[7]  ( .D(
        n12782), .CLK(clk), .Q(
        \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [7]) );
  DFFX1 \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[7]  ( .D(
        \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [7]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [7]) );
  DFFX1 \fadd_0_0_0_0_9/n284_q_reg  ( .D(n12782), .CLK(clk), .Q(
        \fadd_0_0_0_0_9/synceffsub_d1 ) );
  DFFX1 \fadd_0_0_0_0_9/n285_q_reg  ( .D(\fadd_0_0_0_0_9/synceffsub_d1 ), 
        .CLK(clk), .QN(n12095) );
  DFFX1 \fadd_0_0_0_0_9/n276_q_reg  ( .D(n12782), .CLK(clk), .Q(
        \fadd_0_0_0_0_9/effsub_d1 ) );
  DFFX1 \fadd_0_0_0_0_9/n277_q_reg  ( .D(\fadd_0_0_0_0_9/effsub_d1 ), .CLK(clk), .QN(n11596) );
  DFFX1 \p_val_251_reg[11]  ( .D(n12482), .CLK(clk), .Q(n14017) );
  DFFX1 \p_val_296_reg[11]  ( .D(n12481), .CLK(clk), .Q(n14092), .QN(n12097)
         );
  DFFX1 \fadd_0_0_0_0_9_x_reg[11]  ( .D(n12920), .CLK(clk), .Q(n13513), .QN(
        n12784) );
  DFFX1 \fadd_0_0_0_0_9/n293_q_reg[3]  ( .D(\fadd_0_0_0_0_9/newx [11]), .CLK(
        clk), .Q(\fadd_0_0_0_0_9/syncexnxy_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_9/n294_q_reg[3]  ( .D(\fadd_0_0_0_0_9/syncexnxy_d1 [3]), 
        .CLK(clk), .Q(n13776), .QN(n12102) );
  DFFX1 \p_val_251_reg[10]  ( .D(n12480), .CLK(clk), .Q(n14018) );
  DFFX1 \p_val_296_reg[10]  ( .D(n12479), .CLK(clk), .Q(n14093), .QN(n12094)
         );
  DFFX1 \fadd_0_0_0_0_9_x_reg[10]  ( .D(n12921), .CLK(clk), .Q(n13504), .QN(
        n12785) );
  DFFX1 \fadd_0_0_0_0_9/n286_q_reg[9]  ( .D(n14880), .CLK(clk), .Q(
        \fadd_0_0_0_0_9/syncx_d1 [9]) );
  DFFX1 \fadd_0_0_0_0_9/n287_q_reg[9]  ( .D(\fadd_0_0_0_0_9/syncx_d1 [9]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_9/syncx_d2 [9]) );
  DFFX1 \fadd_0_0_0_0_9/n286_q_reg[0]  ( .D(
        \add_0_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .CLK(clk), .Q(\fadd_0_0_0_0_9/syncx_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_9/n287_q_reg[0]  ( .D(\fadd_0_0_0_0_9/syncx_d1 [0]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_9/syncx_d2 [0]) );
  DFFX1 \p_val_251_reg[0]  ( .D(n12478), .CLK(clk), .Q(n14019) );
  DFFX1 \p_val_296_reg[0]  ( .D(n12477), .CLK(clk), .Q(n13793) );
  DFFX1 \fadd_0_0_0_0_9_x_reg[0]  ( .D(n12931), .CLK(clk), .Q(n13521), .QN(
        n11835) );
  DFFX1 \fadd_0_0_0_0_9/rightshiftercomponent/n415_q_reg[2]  ( .D(n14884), 
        .CLK(clk), .QN(n11602) );
  DFFX1 \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/n432_q_reg[2]  ( .D(
        \add_0_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .CLK(clk), .Q(\fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/n433_q_reg[2]  ( .D(
        \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [2]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/x_d2 [2]) );
  DFFX1 \fadd_0_0_0_0_9/n293_q_reg[2]  ( .D(\fadd_0_0_0_0_9/newx [10]), .CLK(
        clk), .Q(\fadd_0_0_0_0_9/syncexnxy_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_9/n294_q_reg[2]  ( .D(\fadd_0_0_0_0_9/syncexnxy_d1 [2]), 
        .CLK(clk), .Q(n13732), .QN(n12100) );
  DFFX1 \fadd_0_0_0_0_9/n286_q_reg[1]  ( .D(
        \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ), .CLK(clk), .Q(\fadd_0_0_0_0_9/syncx_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_9/n287_q_reg[1]  ( .D(\fadd_0_0_0_0_9/syncx_d1 [1]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_9/syncx_d2 [1]) );
  DFFX1 \p_val_251_reg[1]  ( .D(n12476), .CLK(clk), .Q(n14020) );
  DFFX1 \p_val_296_reg[1]  ( .D(n12475), .CLK(clk), .Q(n13794) );
  DFFX1 \fadd_0_0_0_0_9_x_reg[1]  ( .D(n12930), .CLK(clk), .Q(n13532), .QN(
        n11836) );
  DFFX1 \fadd_0_0_0_0_9/rightshiftercomponent/n415_q_reg[3]  ( .D(n14883), 
        .CLK(clk), .QN(n11603) );
  DFFX1 \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/n432_q_reg[3]  ( .D(
        \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ), .CLK(clk), .Q(\fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/n433_q_reg[3]  ( .D(
        \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [3]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/x_d2 [3]) );
  DFFX1 \fadd_0_0_0_0_9/n286_q_reg[2]  ( .D(
        \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ), .CLK(clk), .Q(\fadd_0_0_0_0_9/syncx_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_9/n287_q_reg[2]  ( .D(\fadd_0_0_0_0_9/syncx_d1 [2]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_9/syncx_d2 [2]) );
  DFFX1 \p_val_251_reg[2]  ( .D(n12474), .CLK(clk), .Q(n14021) );
  DFFX1 \p_val_296_reg[2]  ( .D(n12473), .CLK(clk), .Q(n13795) );
  DFFX1 \fadd_0_0_0_0_9_x_reg[2]  ( .D(n12929), .CLK(clk), .Q(n13557), .QN(
        n11837) );
  DFFX1 \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/n432_q_reg[4]  ( .D(
        \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ), .CLK(clk), .Q(\fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/n433_q_reg[4]  ( .D(
        \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [4]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/x_d2 [4]) );
  DFFX1 \fadd_0_0_0_0_9/n286_q_reg[3]  ( .D(
        \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ), .CLK(clk), .Q(\fadd_0_0_0_0_9/syncx_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_9/n287_q_reg[3]  ( .D(\fadd_0_0_0_0_9/syncx_d1 [3]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_9/syncx_d2 [3]) );
  DFFX1 \p_val_251_reg[3]  ( .D(n12472), .CLK(clk), .Q(n14022) );
  DFFX1 \p_val_296_reg[3]  ( .D(n12471), .CLK(clk), .Q(n13796) );
  DFFX1 \fadd_0_0_0_0_9_x_reg[3]  ( .D(n12928), .CLK(clk), .Q(n13574), .QN(
        n11838) );
  DFFX1 \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/n432_q_reg[5]  ( .D(
        \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ), .CLK(clk), .Q(\fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [5]) );
  DFFX1 \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/n433_q_reg[5]  ( .D(
        \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [5]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/x_d2 [5]) );
  DFFX1 \fadd_0_0_0_0_9/n275_q_reg[4]  ( .D(\fadd_0_0_0_0_9/newx [4]), .CLK(
        clk), .Q(\fadd_0_0_0_0_9/newx_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_9/n281_q_reg[0]  ( .D(\fadd_0_0_0_0_9/newx [4]), .CLK(
        clk), .Q(\fadd_0_0_0_0_9/exponentresultfar0_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_9/n282_q_reg[0]  ( .D(
        \fadd_0_0_0_0_9/exponentresultfar0_d1 [0]), .CLK(clk), .Q(
        \fadd_0_0_0_0_9/exponentresultfar0_d2 [0]) );
  DFFX1 \fadd_0_0_0_0_9/n286_q_reg[4]  ( .D(\fadd_0_0_0_0_9/newx [4]), .CLK(
        clk), .Q(\fadd_0_0_0_0_9/syncx_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_9/n287_q_reg[4]  ( .D(\fadd_0_0_0_0_9/syncx_d1 [4]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_9/syncx_d2 [4]) );
  DFFX1 \p_val_251_reg[4]  ( .D(n12470), .CLK(clk), .Q(n14023) );
  DFFX1 \p_val_296_reg[4]  ( .D(n12469), .CLK(clk), .Q(n13797) );
  DFFX1 \fadd_0_0_0_0_9_x_reg[4]  ( .D(n12927), .CLK(clk), .Q(n5346), .QN(
        n14639) );
  DFFX1 \fadd_0_0_0_0_9/n275_q_reg[5]  ( .D(\fadd_0_0_0_0_9/newx [5]), .CLK(
        clk), .Q(\fadd_0_0_0_0_9/newx_d1 [5]) );
  DFFX1 \fadd_0_0_0_0_9/n281_q_reg[1]  ( .D(\fadd_0_0_0_0_9/newx [5]), .CLK(
        clk), .Q(\fadd_0_0_0_0_9/exponentresultfar0_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_9/n282_q_reg[1]  ( .D(
        \fadd_0_0_0_0_9/exponentresultfar0_d1 [1]), .CLK(clk), .Q(
        \fadd_0_0_0_0_9/exponentresultfar0_d2 [1]) );
  DFFX1 \fadd_0_0_0_0_9/n286_q_reg[5]  ( .D(\fadd_0_0_0_0_9/newx [5]), .CLK(
        clk), .Q(\fadd_0_0_0_0_9/syncx_d1 [5]) );
  DFFX1 \fadd_0_0_0_0_9/n287_q_reg[5]  ( .D(\fadd_0_0_0_0_9/syncx_d1 [5]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_9/syncx_d2 [5]) );
  DFFX1 \p_val_251_reg[5]  ( .D(n12468), .CLK(clk), .Q(n14024) );
  DFFX1 \p_val_296_reg[5]  ( .D(n12467), .CLK(clk), .Q(n13798) );
  DFFX1 \fadd_0_0_0_0_9_x_reg[5]  ( .D(n12926), .CLK(clk), .Q(n5347), .QN(
        n14638) );
  DFFX1 \fadd_0_0_0_0_9/n275_q_reg[6]  ( .D(\fadd_0_0_0_0_9/newx [6]), .CLK(
        clk), .Q(\fadd_0_0_0_0_9/newx_d1 [6]) );
  DFFX1 \fadd_0_0_0_0_9/n281_q_reg[2]  ( .D(\fadd_0_0_0_0_9/newx [6]), .CLK(
        clk), .Q(\fadd_0_0_0_0_9/exponentresultfar0_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_9/n282_q_reg[2]  ( .D(
        \fadd_0_0_0_0_9/exponentresultfar0_d1 [2]), .CLK(clk), .Q(
        \fadd_0_0_0_0_9/exponentresultfar0_d2 [2]) );
  DFFX1 \fadd_0_0_0_0_9/n286_q_reg[6]  ( .D(\fadd_0_0_0_0_9/newx [6]), .CLK(
        clk), .Q(\fadd_0_0_0_0_9/syncx_d1 [6]) );
  DFFX1 \fadd_0_0_0_0_9/n287_q_reg[6]  ( .D(\fadd_0_0_0_0_9/syncx_d1 [6]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_9/syncx_d2 [6]) );
  DFFX1 \p_val_251_reg[6]  ( .D(n12466), .CLK(clk), .Q(n14025) );
  DFFX1 \p_val_296_reg[6]  ( .D(n12465), .CLK(clk), .Q(n13799) );
  DFFX1 \fadd_0_0_0_0_9_x_reg[6]  ( .D(n12925), .CLK(clk), .Q(n5348), .QN(
        n14637) );
  DFFX1 \fadd_0_0_0_0_9/n275_q_reg[7]  ( .D(\fadd_0_0_0_0_9/newx [7]), .CLK(
        clk), .Q(\fadd_0_0_0_0_9/newx_d1 [7]) );
  DFFX1 \fadd_0_0_0_0_9/n281_q_reg[3]  ( .D(\fadd_0_0_0_0_9/newx [7]), .CLK(
        clk), .Q(\fadd_0_0_0_0_9/exponentresultfar0_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_9/n282_q_reg[3]  ( .D(
        \fadd_0_0_0_0_9/exponentresultfar0_d1 [3]), .CLK(clk), .Q(
        \fadd_0_0_0_0_9/exponentresultfar0_d2 [3]) );
  DFFX1 \fadd_0_0_0_0_9/n286_q_reg[7]  ( .D(\fadd_0_0_0_0_9/newx [7]), .CLK(
        clk), .Q(\fadd_0_0_0_0_9/syncx_d1 [7]) );
  DFFX1 \fadd_0_0_0_0_9/n287_q_reg[7]  ( .D(\fadd_0_0_0_0_9/syncx_d1 [7]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_9/syncx_d2 [7]) );
  DFFX1 \p_val_251_reg[7]  ( .D(n12464), .CLK(clk), .Q(n14026) );
  DFFX1 \p_val_296_reg[7]  ( .D(n12463), .CLK(clk), .Q(n13800) );
  DFFX1 \fadd_0_0_0_0_9_x_reg[7]  ( .D(n12924), .CLK(clk), .Q(n5349), .QN(
        n14636) );
  DFFX1 \fadd_0_0_0_0_9/n275_q_reg[8]  ( .D(\fadd_0_0_0_0_9/newx [8]), .CLK(
        clk), .Q(\fadd_0_0_0_0_9/newx_d1 [8]) );
  DFFX1 \fadd_0_0_0_0_9/n280_q_reg[0]  ( .D(
        \fadd_0_0_0_0_9/exponentresultclose [0]), .CLK(clk), .Q(
        \fadd_0_0_0_0_9/exponentresultclose_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_9/n280_q_reg[1]  ( .D(
        \fadd_0_0_0_0_9/exponentresultclose [1]), .CLK(clk), .Q(
        \fadd_0_0_0_0_9/exponentresultclose_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_9/n280_q_reg[2]  ( .D(
        \fadd_0_0_0_0_9/exponentresultclose [2]), .CLK(clk), .Q(
        \fadd_0_0_0_0_9/exponentresultclose_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_9/n280_q_reg[3]  ( .D(
        \fadd_0_0_0_0_9/exponentresultclose [3]), .CLK(clk), .Q(
        \fadd_0_0_0_0_9/exponentresultclose_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_9/n280_q_reg[4]  ( .D(
        \fadd_0_0_0_0_9/exponentresultclose [4]), .CLK(clk), .Q(
        \fadd_0_0_0_0_9/exponentresultclose_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_9/n280_q_reg[6]  ( .D(n13655), .CLK(clk), .Q(
        \fadd_0_0_0_0_9/exponentresultclose_d1 [6]) );
  DFFX1 \fadd_0_0_0_0_9/n280_q_reg[5]  ( .D(n13655), .CLK(clk), .Q(
        \fadd_0_0_0_0_9/exponentresultclose_d1 [5]) );
  DFFX1 \fadd_0_0_0_0_9/n281_q_reg[4]  ( .D(\fadd_0_0_0_0_9/newx [8]), .CLK(
        clk), .Q(\fadd_0_0_0_0_9/exponentresultfar0_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_9/n282_q_reg[4]  ( .D(
        \fadd_0_0_0_0_9/exponentresultfar0_d1 [4]), .CLK(clk), .Q(
        \fadd_0_0_0_0_9/exponentresultfar0_d2 [4]) );
  DFFX1 \fadd_0_0_0_0_9/n286_q_reg[8]  ( .D(\fadd_0_0_0_0_9/newx [8]), .CLK(
        clk), .Q(\fadd_0_0_0_0_9/syncx_d1 [8]) );
  DFFX1 \fadd_0_0_0_0_9/n287_q_reg[8]  ( .D(\fadd_0_0_0_0_9/syncx_d1 [8]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_9/syncx_d2 [8]) );
  DFFX1 \p_val_251_reg[8]  ( .D(n12462), .CLK(clk), .Q(n14027) );
  DFFX1 \p_val_296_reg[8]  ( .D(n12461), .CLK(clk), .Q(n13801) );
  DFFX1 \fadd_0_0_0_0_9_x_reg[8]  ( .D(n12923), .CLK(clk), .Q(n5350), .QN(
        n14635) );
  DFFX1 \fadd_0_0_0_0_9/rightshiftercomponent/n413_q_reg[2]  ( .D(n14874), 
        .CLK(clk), .Q(\fadd_0_0_0_0_9/rightshiftercomponent/ps_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_9/rightshiftercomponent/n416_q_reg[1]  ( .D(
        \fadd_0_0_0_0_9/rightshiftercomponent/level2[1] ), .CLK(clk), .QN(
        n11604) );
  DFFX1 \fadd_0_0_0_0_9/rightshiftercomponent/n416_q_reg[0]  ( .D(n12781), 
        .CLK(clk), .QN(n11605) );
  DFFX1 \fadd_0_0_0_0_9/rightshiftercomponent/n413_q_reg[1]  ( .D(n14877), 
        .CLK(clk), .Q(\fadd_0_0_0_0_9/rightshiftercomponent/ps_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_9/rightshiftercomponent/n417_q_reg  ( .D(
        \fadd_0_0_0_0_9/rightshiftercomponent/n389_o ), .CLK(clk), .Q(n14960)
         );
  DFFX1 \fadd_0_0_0_0_9/rightshiftercomponent/n418_q_reg[0]  ( .D(n12780), 
        .CLK(clk), .Q(\fadd_0_0_0_0_9/rightshiftercomponent/level1_d1[0] ) );
  DFFX1 \fadd_0_0_0_0_9/rightshiftercomponent/n419_q_reg[0]  ( .D(
        \fadd_0_0_0_0_9/rightshiftercomponent/level1_d1[0] ), .CLK(clk), .Q(
        \fadd_0_0_0_0_9/rightshiftercomponent/level1_d2[0] ) );
  DFFX1 \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[5]  ( .D(
        \fadd_0_0_0_0_9/fracyfarxorop [5]), .CLK(clk), .Q(
        \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [5]) );
  DFFX1 \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[5]  ( .D(
        \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [5]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [5]) );
  DFFX1 \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[3]  ( .D(
        \fadd_0_0_0_0_9/fracyfarxorop [3]), .CLK(clk), .Q(
        \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[3]  ( .D(
        \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [3]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [3]) );
  DFFX1 \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[2]  ( .D(
        \fadd_0_0_0_0_9/fracyfarxorop [2]), .CLK(clk), .Q(
        \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[2]  ( .D(
        \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [2]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [2]) );
  DFFX1 \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[1]  ( .D(
        \fadd_0_0_0_0_9/fracyfarxorop [1]), .CLK(clk), .Q(
        \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[1]  ( .D(
        \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [1]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [1]) );
  DFFX1 \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[0]  ( .D(
        \fadd_0_0_0_0_9/fracyfarxorop [0]), .CLK(clk), .Q(
        \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[0]  ( .D(
        \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [0]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [0]) );
  DFFX1 \fadd_0_0_0_0_9/rightshiftercomponent/n413_q_reg[0]  ( .D(n12779), 
        .CLK(clk), .Q(\fadd_0_0_0_0_9/rightshiftercomponent/ps_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_9/rightshiftercomponent/n414_q_reg[0]  ( .D(
        \fadd_0_0_0_0_9/rightshiftercomponent/ps_d1 [0]), .CLK(clk), .Q(
        \fadd_0_0_0_0_9/rightshiftercomponent/ps_d2[0] ) );
  DFFX1 \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[4]  ( .D(
        \fadd_0_0_0_0_9/fracyfarxorop [4]), .CLK(clk), .Q(
        \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[4]  ( .D(
        \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [4]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [4]) );
  DFFX1 \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[6]  ( .D(
        \fadd_0_0_0_0_9/fracyfarxorop [6]), .CLK(clk), .Q(
        \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [6]) );
  DFFX1 \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[6]  ( .D(
        \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [6]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [6]) );
  DFFX1 \fadd_0_0_0_0_9/n293_q_reg[1]  ( .D(\fadd_0_0_0_0_9/newy_11 ), .CLK(
        clk), .Q(\fadd_0_0_0_0_9/syncexnxy_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_9/n294_q_reg[1]  ( .D(\fadd_0_0_0_0_9/syncexnxy_d1 [1]), 
        .CLK(clk), .Q(n13739), .QN(n12103) );
  DFFX1 \fadd_0_0_0_0_9/n278_q_reg  ( .D(n14873), .CLK(clk), .Q(
        \fadd_0_0_0_0_9/selectclosepath_d1 ), .QN(n11607) );
  DFFX1 \fadd_0_0_0_0_9/n283_q_reg  ( .D(\fadd_0_0_0_0_9/zerofromclose ), 
        .CLK(clk), .Q(\fadd_0_0_0_0_9/zerofromclose_d1 ) );
  DFFX1 \fadd_0_0_0_0_9/n290_q_reg  ( .D(\fadd_0_0_0_0_9/ressign ), .CLK(clk), 
        .Q(\fadd_0_0_0_0_9/syncressign_d1 ) );
  DFFX1 \fadd_0_0_0_0_9/n291_q_reg  ( .D(\fadd_0_0_0_0_9/syncressign_d1 ), 
        .CLK(clk), .QN(n12105) );
  DFFX1 \fmul_0_0_0_0_10/roundingadder/n155_q_reg[0]  ( .D(
        \fmul_0_0_0_0_10/U8/Z_5 ), .CLK(clk), .Q(
        \fmul_0_0_0_0_10/roundingadder/add_1_root_add_57/A[0] ) );
  DFFX1 \fmul_0_0_0_0_10/roundingadder/n155_q_reg[1]  ( .D(
        \fmul_0_0_0_0_10/U8/Z_6 ), .CLK(clk), .Q(
        \fmul_0_0_0_0_10/roundingadder/add_1_root_add_57/A[1] ) );
  DFFX1 \fmul_0_0_0_0_10/roundingadder/n155_q_reg[2]  ( .D(
        \fmul_0_0_0_0_10/U8/Z_7 ), .CLK(clk), .Q(
        \fmul_0_0_0_0_10/roundingadder/add_1_root_add_57/A[2] ) );
  DFFX1 \fmul_0_0_0_0_10/roundingadder/n155_q_reg[3]  ( .D(
        \fmul_0_0_0_0_10/U8/Z_8 ), .CLK(clk), .Q(
        \fmul_0_0_0_0_10/roundingadder/add_1_root_add_57/A[3] ) );
  DFFX1 \fmul_0_0_0_0_10/roundingadder/n155_q_reg[4]  ( .D(n14919), .CLK(clk), 
        .Q(\fmul_0_0_0_0_10/roundingadder/add_1_root_add_57/A[4] ) );
  DFFX1 \fmul_0_0_0_0_10/roundingadder/n155_q_reg[5]  ( .D(
        \fmul_0_0_0_0_10/sub_1_root_add_321/DIFF[1] ), .CLK(clk), .Q(
        \fmul_0_0_0_0_10/roundingadder/add_1_root_add_57/A[5] ) );
  DFFX1 \fmul_0_0_0_0_10/roundingadder/n155_q_reg[6]  ( .D(
        \fmul_0_0_0_0_10/sub_1_root_add_321/DIFF[2] ), .CLK(clk), .Q(
        \fmul_0_0_0_0_10/roundingadder/add_1_root_add_57/A[6] ) );
  DFFX1 \fmul_0_0_0_0_10/roundingadder/n155_q_reg[7]  ( .D(
        \fmul_0_0_0_0_10/sub_1_root_add_321/DIFF[3] ), .CLK(clk), .Q(
        \fmul_0_0_0_0_10/roundingadder/add_1_root_add_57/A[7] ) );
  DFFX1 \fmul_0_0_0_0_10/roundingadder/n155_q_reg[8]  ( .D(
        \fmul_0_0_0_0_10/sub_1_root_add_321/DIFF[4] ), .CLK(clk), .Q(
        \fmul_0_0_0_0_10/roundingadder/add_1_root_add_57/A[8] ) );
  DFFX1 \fmul_0_0_0_0_10/roundingadder/n155_q_reg[9]  ( .D(
        \fmul_0_0_0_0_10/sub_1_root_add_321/DIFF[5] ), .CLK(clk), .Q(
        \fmul_0_0_0_0_10/roundingadder/add_1_root_add_57/A[9] ) );
  DFFX1 \fmul_0_0_0_0_10/roundingadder/n155_q_reg[10]  ( .D(n14119), .CLK(clk), 
        .QN(n14150) );
  DFFX1 \fmul_0_0_0_0_10/roundingadder/n154_q_reg  ( .D(\fmul_0_0_0_0_10/n98 ), 
        .CLK(clk), .Q(\fmul_0_0_0_0_10/roundingadder/add_1_root_add_57/CI ) );
  DFFX1 \fadd_0_0_0_0_10_y_reg[0]  ( .D(n12919), .CLK(clk), .Q(n13633), .QN(
        n11845) );
  DFFX1 \fadd_0_0_0_0_10_y_reg[1]  ( .D(n12918), .CLK(clk), .Q(n13646), .QN(
        n11846) );
  DFFX1 \fadd_0_0_0_0_10_y_reg[2]  ( .D(n12917), .CLK(clk), .Q(n13673), .QN(
        n11847) );
  DFFX1 \fadd_0_0_0_0_10_y_reg[3]  ( .D(n12916), .CLK(clk), .Q(n13696), .QN(
        n11848) );
  DFFX1 \fadd_0_0_0_0_10_y_reg[4]  ( .D(n12915), .CLK(clk), .Q(n13885), .QN(
        n14179) );
  DFFX1 \fadd_0_0_0_0_10_y_reg[5]  ( .D(n12914), .CLK(clk), .Q(n14980), .QN(
        n12813) );
  DFFX1 \fadd_0_0_0_0_10_y_reg[6]  ( .D(n12913), .CLK(clk), .Q(n14981), .QN(
        n12812) );
  DFFX1 \fadd_0_0_0_0_10_y_reg[7]  ( .D(n12912), .CLK(clk), .Q(n14982), .QN(
        n12811) );
  DFFX1 \fadd_0_0_0_0_10_y_reg[8]  ( .D(n12911), .CLK(clk), .Q(n14983), .QN(
        n12810) );
  DFFX1 \fadd_0_0_0_0_10_y_reg[11]  ( .D(n12908), .CLK(clk), .Q(n13886), .QN(
        n12808) );
  DFFX1 \fadd_0_0_0_0_10_y_reg[10]  ( .D(n12909), .CLK(clk), .Q(n13887), .QN(
        n12809) );
  DFFX1 \fadd_0_0_0_0_10/n286_q_reg[8]  ( .D(\fadd_0_0_0_0_10/U29/Z_8 ), .CLK(
        clk), .Q(\fadd_0_0_0_0_10/n167 ) );
  DFFX1 \fadd_0_0_0_0_10/n287_q_reg[8]  ( .D(\fadd_0_0_0_0_10/n167 ), .CLK(clk), .Q(\fadd_0_0_0_0_10/U11/DATA2_8 ) );
  DFFX1 \fadd_0_0_0_0_10/n281_q_reg[4]  ( .D(\fadd_0_0_0_0_10/U29/Z_8 ), .CLK(
        clk), .Q(\fadd_0_0_0_0_10/n213 ) );
  DFFX1 \fadd_0_0_0_0_10/n282_q_reg[4]  ( .D(\fadd_0_0_0_0_10/n213 ), .CLK(clk), .QN(n12067) );
  DFFX1 \fadd_0_0_0_0_10/n275_q_reg[8]  ( .D(\fadd_0_0_0_0_10/U29/Z_8 ), .CLK(
        clk), .QN(n13884) );
  DFFX1 \fadd_0_0_0_0_10/n280_q_reg[4]  ( .D(\fadd_0_0_0_0_10/sub_784/DIFF[4] ), .CLK(clk), .QN(n12024) );
  DFFX1 \fadd_0_0_0_0_10/n280_q_reg[5]  ( .D(n14126), .CLK(clk), .Q(
        \fadd_0_0_0_0_10/U4/DATA1_9 ) );
  DFFX1 \fadd_0_0_0_0_10/n280_q_reg[6]  ( .D(n14126), .CLK(clk), .Q(
        \fadd_0_0_0_0_10/U4/DATA1_10 ) );
  DFFX1 \p_val_275_reg[10]  ( .D(n12460), .CLK(clk), .Q(n14028) );
  DFFX1 \p_val_297_reg[10]  ( .D(n12459), .CLK(clk), .Q(n14078), .QN(n12066)
         );
  DFFX1 \p_val_307_reg[10]  ( .D(n12458), .CLK(clk), .QN(n12065) );
  DFFX1 \fadd_0_0_0_0_10_x_reg[10]  ( .D(n12897), .CLK(clk), .Q(n13469) );
  DFFX1 \fadd_0_0_0_0_10/n293_q_reg[0]  ( .D(\fadd_0_0_0_0_10/U28/Z_5 ), .CLK(
        clk), .Q(\fadd_0_0_0_0_10/n142 ) );
  DFFX1 \fadd_0_0_0_0_10/n294_q_reg[0]  ( .D(\fadd_0_0_0_0_10/n142 ), .CLK(clk), .Q(n12073), .QN(n13745) );
  DFFX1 \fadd_0_0_0_0_10/n293_q_reg[2]  ( .D(\fadd_0_0_0_0_10/U29/Z_10 ), 
        .CLK(clk), .Q(\fadd_0_0_0_0_10/n144 ) );
  DFFX1 \fadd_0_0_0_0_10/n294_q_reg[2]  ( .D(\fadd_0_0_0_0_10/n144 ), .CLK(clk), .Q(n13724) );
  DFFX1 \p_val_275_reg[0]  ( .D(n12457), .CLK(clk), .Q(n14029) );
  DFFX1 \p_val_297_reg[0]  ( .D(n12456), .CLK(clk), .Q(n14058) );
  DFFX1 \p_val_307_reg[0]  ( .D(n12455), .CLK(clk), .Q(n13596) );
  DFFX1 \fadd_0_0_0_0_10_x_reg[0]  ( .D(n12907), .CLK(clk), .Q(n13477), .QN(
        n11850) );
  DFFX1 \fadd_0_0_0_0_10/rightshiftercomponent/n415_q_reg[2]  ( .D(n14965), 
        .CLK(clk), .QN(n11500) );
  DFFX1 \fadd_0_0_0_0_10/n286_q_reg[0]  ( .D(\fadd_0_0_0_0_10/U29/Z_0 ), .CLK(
        clk), .Q(\fadd_0_0_0_0_10/n159 ) );
  DFFX1 \fadd_0_0_0_0_10/n287_q_reg[0]  ( .D(\fadd_0_0_0_0_10/n159 ), .CLK(clk), .Q(\fadd_0_0_0_0_10/U11/DATA2_0 ) );
  DFFX1 \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/n432_q_reg[2]  ( .D(
        \fadd_0_0_0_0_10/U29/Z_0 ), .CLK(clk), .Q(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/n433_q_reg[2]  ( .D(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [2]), .CLK(clk), 
        .Q(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/A[2] ) );
  DFFX1 \fadd_0_0_0_0_10/norm/n351_q_reg[5]  ( .D(\fadd_0_0_0_0_10/U24/Z_5 ), 
        .CLK(clk), .QN(n11887) );
  DFFX1 \fadd_0_0_0_0_10/n290_q_reg  ( .D(\fadd_0_0_0_0_10/U23/Z_0 ), .CLK(clk), .Q(\fadd_0_0_0_0_10/n146 ) );
  DFFX1 \fadd_0_0_0_0_10/n291_q_reg  ( .D(\fadd_0_0_0_0_10/n146 ), .CLK(clk), 
        .QN(n12057) );
  DFFX1 \p_val_275_reg[9]  ( .D(n12454), .CLK(clk), .Q(n14030) );
  DFFX1 \p_val_297_reg[9]  ( .D(n12453), .CLK(clk), .Q(n14079), .QN(n12056) );
  DFFX1 \p_val_307_reg[9]  ( .D(n12452), .CLK(clk), .QN(n12055) );
  DFFX1 \fadd_0_0_0_0_10_x_reg[9]  ( .D(n12898), .CLK(clk), .Q(n13585), .QN(
        n11854) );
  DFFX1 \fadd_0_0_0_0_10/n288_q_reg  ( .D(\fadd_0_0_0_0_10/U28/Z_4 ), .CLK(clk), .Q(\fadd_0_0_0_0_10/n148 ) );
  DFFX1 \fadd_0_0_0_0_10/n289_q_reg  ( .D(\fadd_0_0_0_0_10/n148 ), .CLK(clk), 
        .Q(\fadd_0_0_0_0_10/n147 ) );
  DFFX1 \fadd_0_0_0_0_10/n286_q_reg[9]  ( .D(n14940), .CLK(clk), .Q(
        \fadd_0_0_0_0_10/n168 ) );
  DFFX1 \fadd_0_0_0_0_10/n287_q_reg[9]  ( .D(\fadd_0_0_0_0_10/n168 ), .CLK(clk), .Q(\fadd_0_0_0_0_10/U12/DATA3_0 ) );
  DFFX1 \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[7]  ( .D(
        n14938), .CLK(clk), .Q(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [7]) );
  DFFX1 \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[7]  ( .D(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [7]), .CLK(clk), 
        .Q(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/B[7] ) );
  DFFX1 \fadd_0_0_0_0_10/n276_q_reg  ( .D(n14938), .CLK(clk), .Q(
        \fadd_0_0_0_0_10/n305 ) );
  DFFX1 \fadd_0_0_0_0_10/n277_q_reg  ( .D(\fadd_0_0_0_0_10/n305 ), .CLK(clk), 
        .QN(n11496) );
  DFFX1 \p_val_275_reg[1]  ( .D(n12451), .CLK(clk), .Q(n14031) );
  DFFX1 \p_val_297_reg[1]  ( .D(n12450), .CLK(clk), .Q(n14059) );
  DFFX1 \p_val_307_reg[1]  ( .D(n12449), .CLK(clk), .Q(n13597) );
  DFFX1 \fadd_0_0_0_0_10_x_reg[1]  ( .D(n12906), .CLK(clk), .Q(n13526), .QN(
        n11851) );
  DFFX1 \fadd_0_0_0_0_10/rightshiftercomponent/n415_q_reg[3]  ( .D(n14968), 
        .CLK(clk), .QN(n11501) );
  DFFX1 \fadd_0_0_0_0_10/n286_q_reg[1]  ( .D(\fadd_0_0_0_0_10/U29/Z_1 ), .CLK(
        clk), .Q(\fadd_0_0_0_0_10/n160 ) );
  DFFX1 \fadd_0_0_0_0_10/n287_q_reg[1]  ( .D(\fadd_0_0_0_0_10/n160 ), .CLK(clk), .Q(\fadd_0_0_0_0_10/U11/DATA2_1 ) );
  DFFX1 \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/n432_q_reg[3]  ( .D(
        \fadd_0_0_0_0_10/U29/Z_1 ), .CLK(clk), .Q(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/n433_q_reg[3]  ( .D(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [3]), .CLK(clk), 
        .Q(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/A[3] ) );
  DFFX1 \p_val_275_reg[2]  ( .D(n12448), .CLK(clk), .Q(n14032) );
  DFFX1 \p_val_297_reg[2]  ( .D(n12447), .CLK(clk), .Q(n14060) );
  DFFX1 \p_val_307_reg[2]  ( .D(n12446), .CLK(clk), .Q(n13598) );
  DFFX1 \fadd_0_0_0_0_10_x_reg[2]  ( .D(n12905), .CLK(clk), .Q(n13538), .QN(
        n11852) );
  DFFX1 \fadd_0_0_0_0_10/n286_q_reg[2]  ( .D(\fadd_0_0_0_0_10/U29/Z_2 ), .CLK(
        clk), .Q(\fadd_0_0_0_0_10/n161 ) );
  DFFX1 \fadd_0_0_0_0_10/n287_q_reg[2]  ( .D(\fadd_0_0_0_0_10/n161 ), .CLK(clk), .Q(\fadd_0_0_0_0_10/U11/DATA2_2 ) );
  DFFX1 \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/n432_q_reg[4]  ( .D(
        \fadd_0_0_0_0_10/U29/Z_2 ), .CLK(clk), .Q(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/n433_q_reg[4]  ( .D(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [4]), .CLK(clk), 
        .Q(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/A[4] ) );
  DFFX1 \p_val_275_reg[3]  ( .D(n12445), .CLK(clk), .Q(n14033) );
  DFFX1 \p_val_297_reg[3]  ( .D(n12444), .CLK(clk), .Q(n14061) );
  DFFX1 \p_val_307_reg[3]  ( .D(n12443), .CLK(clk), .Q(n13599) );
  DFFX1 \fadd_0_0_0_0_10_x_reg[3]  ( .D(n12904), .CLK(clk), .Q(n13562), .QN(
        n11853) );
  DFFX1 \fadd_0_0_0_0_10/n286_q_reg[3]  ( .D(\fadd_0_0_0_0_10/U29/Z_3 ), .CLK(
        clk), .Q(\fadd_0_0_0_0_10/n162 ) );
  DFFX1 \fadd_0_0_0_0_10/n287_q_reg[3]  ( .D(\fadd_0_0_0_0_10/n162 ), .CLK(clk), .Q(\fadd_0_0_0_0_10/U11/DATA2_3 ) );
  DFFX1 \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/n432_q_reg[5]  ( .D(
        \fadd_0_0_0_0_10/U29/Z_3 ), .CLK(clk), .Q(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [5]) );
  DFFX1 \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/n433_q_reg[5]  ( .D(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [5]), .CLK(clk), 
        .Q(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/A[5] ) );
  DFFX1 \p_val_275_reg[4]  ( .D(n12442), .CLK(clk), .Q(n14034) );
  DFFX1 \p_val_297_reg[4]  ( .D(n12441), .CLK(clk), .Q(n14062) );
  DFFX1 \p_val_307_reg[4]  ( .D(n12440), .CLK(clk), .Q(n13600) );
  DFFX1 \fadd_0_0_0_0_10_x_reg[4]  ( .D(n12903), .CLK(clk), .Q(n13635), .QN(
        n14180) );
  DFFX1 \fadd_0_0_0_0_10/n286_q_reg[4]  ( .D(\fadd_0_0_0_0_10/U29/Z_4 ), .CLK(
        clk), .Q(\fadd_0_0_0_0_10/n163 ) );
  DFFX1 \fadd_0_0_0_0_10/n287_q_reg[4]  ( .D(\fadd_0_0_0_0_10/n163 ), .CLK(clk), .QN(n12042) );
  DFFX1 \fadd_0_0_0_0_10/n281_q_reg[0]  ( .D(\fadd_0_0_0_0_10/U29/Z_4 ), .CLK(
        clk), .Q(\fadd_0_0_0_0_10/n209 ) );
  DFFX1 \fadd_0_0_0_0_10/n282_q_reg[0]  ( .D(\fadd_0_0_0_0_10/n209 ), .CLK(clk), .Q(n13697), .QN(n12041) );
  DFFX1 \fadd_0_0_0_0_10/n275_q_reg[4]  ( .D(\fadd_0_0_0_0_10/U29/Z_4 ), .CLK(
        clk), .QN(n13714) );
  DFFX1 \fadd_0_0_0_0_10/norm/n351_q_reg[2]  ( .D(\fadd_0_0_0_0_10/U24/Z_2 ), 
        .CLK(clk), .QN(n11890) );
  DFFX1 \fadd_0_0_0_0_10/norm/n351_q_reg[3]  ( .D(\fadd_0_0_0_0_10/U24/Z_3 ), 
        .CLK(clk), .QN(n11889) );
  DFFX1 \fadd_0_0_0_0_10/norm/n351_q_reg[4]  ( .D(\fadd_0_0_0_0_10/U24/Z_4 ), 
        .CLK(clk), .QN(n11888) );
  DFFX1 \fadd_0_0_0_0_10/norm/n351_q_reg[1]  ( .D(\fadd_0_0_0_0_10/U24/Z_1 ), 
        .CLK(clk), .QN(n11499) );
  DFFX1 \fadd_0_0_0_0_10/norm/n351_q_reg[0]  ( .D(n14964), .CLK(clk), .QN(
        n11498) );
  DFFX1 \fadd_0_0_0_0_10/n280_q_reg[0]  ( .D(\fadd_0_0_0_0_10/sub_784/DIFF[0] ), .CLK(clk), .Q(\fadd_0_0_0_0_10/U4/DATA1_4 ) );
  DFFX1 \fadd_0_0_0_0_10/norm/n353_q_reg  ( .D(n14178), .CLK(clk), .QN(n12061)
         );
  DFFX1 \fadd_0_0_0_0_10/norm/n352_q_reg[4]  ( .D(
        \fadd_0_0_0_0_10/norm/U5/Z_4 ), .CLK(clk), .Q(
        \fadd_0_0_0_0_10/norm/U4/DATA2_5 ) );
  DFFX1 \fadd_0_0_0_0_10/norm/n352_q_reg[3]  ( .D(
        \fadd_0_0_0_0_10/norm/U5/Z_3 ), .CLK(clk), .Q(n13695) );
  DFFX1 \fadd_0_0_0_0_10/norm/n352_q_reg[1]  ( .D(
        \fadd_0_0_0_0_10/norm/U5/Z_1 ), .CLK(clk), .Q(n13485), .QN(n12063) );
  DFFX1 \fadd_0_0_0_0_10/norm/n352_q_reg[0]  ( .D(
        \fadd_0_0_0_0_10/norm/U5/Z_0 ), .CLK(clk), .Q(n13676), .QN(n12062) );
  DFFX1 \fadd_0_0_0_0_10/norm/n352_q_reg[2]  ( .D(
        \fadd_0_0_0_0_10/norm/U5/Z_2 ), .CLK(clk), .Q(n13549) );
  DFFX1 \p_val_275_reg[5]  ( .D(n12439), .CLK(clk), .Q(n14035) );
  DFFX1 \p_val_297_reg[5]  ( .D(n12438), .CLK(clk), .Q(n14063) );
  DFFX1 \p_val_307_reg[5]  ( .D(n12437), .CLK(clk), .Q(n13601) );
  DFFX1 \fadd_0_0_0_0_10_x_reg[5]  ( .D(n12902), .CLK(clk), .Q(n14996), .QN(
        n12806) );
  DFFX1 \fadd_0_0_0_0_10/n286_q_reg[5]  ( .D(\fadd_0_0_0_0_10/U29/Z_5 ), .CLK(
        clk), .Q(\fadd_0_0_0_0_10/n164 ) );
  DFFX1 \fadd_0_0_0_0_10/n287_q_reg[5]  ( .D(\fadd_0_0_0_0_10/n164 ), .CLK(clk), .Q(\fadd_0_0_0_0_10/U11/DATA2_5 ) );
  DFFX1 \fadd_0_0_0_0_10/n281_q_reg[1]  ( .D(\fadd_0_0_0_0_10/U29/Z_5 ), .CLK(
        clk), .Q(\fadd_0_0_0_0_10/n210 ) );
  DFFX1 \fadd_0_0_0_0_10/n282_q_reg[1]  ( .D(\fadd_0_0_0_0_10/n210 ), .CLK(clk), .Q(n13677), .QN(n12036) );
  DFFX1 \fadd_0_0_0_0_10/n275_q_reg[5]  ( .D(\fadd_0_0_0_0_10/U29/Z_5 ), .CLK(
        clk), .Q(\fadd_0_0_0_0_10/sub_784/A[1] ) );
  DFFX1 \fadd_0_0_0_0_10/n280_q_reg[1]  ( .D(\fadd_0_0_0_0_10/sub_784/DIFF[1] ), .CLK(clk), .QN(n12037) );
  DFFX1 \p_val_275_reg[6]  ( .D(n12436), .CLK(clk), .Q(n14036) );
  DFFX1 \p_val_297_reg[6]  ( .D(n12435), .CLK(clk), .Q(n14064) );
  DFFX1 \p_val_307_reg[6]  ( .D(n12434), .CLK(clk), .Q(n13602) );
  DFFX1 \fadd_0_0_0_0_10_x_reg[6]  ( .D(n12901), .CLK(clk), .Q(n14997), .QN(
        n12805) );
  DFFX1 \fadd_0_0_0_0_10/n286_q_reg[6]  ( .D(\fadd_0_0_0_0_10/U29/Z_6 ), .CLK(
        clk), .Q(\fadd_0_0_0_0_10/n165 ) );
  DFFX1 \fadd_0_0_0_0_10/n287_q_reg[6]  ( .D(\fadd_0_0_0_0_10/n165 ), .CLK(clk), .Q(\fadd_0_0_0_0_10/U11/DATA2_6 ) );
  DFFX1 \fadd_0_0_0_0_10/n281_q_reg[2]  ( .D(\fadd_0_0_0_0_10/U29/Z_6 ), .CLK(
        clk), .Q(\fadd_0_0_0_0_10/n211 ) );
  DFFX1 \fadd_0_0_0_0_10/n282_q_reg[2]  ( .D(\fadd_0_0_0_0_10/n211 ), .CLK(clk), .Q(n13706), .QN(n12032) );
  DFFX1 \fadd_0_0_0_0_10/n275_q_reg[6]  ( .D(\fadd_0_0_0_0_10/U29/Z_6 ), .CLK(
        clk), .Q(\fadd_0_0_0_0_10/sub_784/A[2] ) );
  DFFX1 \fadd_0_0_0_0_10/n280_q_reg[2]  ( .D(\fadd_0_0_0_0_10/sub_784/DIFF[2] ), .CLK(clk), .Q(\fadd_0_0_0_0_10/U4/DATA1_6 ) );
  DFFX1 \p_val_275_reg[7]  ( .D(n12433), .CLK(clk), .Q(n14037) );
  DFFX1 \p_val_297_reg[7]  ( .D(n12432), .CLK(clk), .Q(n14065) );
  DFFX1 \p_val_307_reg[7]  ( .D(n12431), .CLK(clk), .Q(n13603) );
  DFFX1 \fadd_0_0_0_0_10_x_reg[7]  ( .D(n12900), .CLK(clk), .Q(n14998), .QN(
        n12804) );
  DFFX1 \fadd_0_0_0_0_10/n286_q_reg[7]  ( .D(\fadd_0_0_0_0_10/U29/Z_7 ), .CLK(
        clk), .Q(\fadd_0_0_0_0_10/n166 ) );
  DFFX1 \fadd_0_0_0_0_10/n287_q_reg[7]  ( .D(\fadd_0_0_0_0_10/n166 ), .CLK(clk), .Q(\fadd_0_0_0_0_10/U11/DATA2_7 ) );
  DFFX1 \fadd_0_0_0_0_10/n281_q_reg[3]  ( .D(\fadd_0_0_0_0_10/U29/Z_7 ), .CLK(
        clk), .Q(\fadd_0_0_0_0_10/n212 ) );
  DFFX1 \fadd_0_0_0_0_10/n282_q_reg[3]  ( .D(\fadd_0_0_0_0_10/n212 ), .CLK(clk), .Q(n13722), .QN(n12028) );
  DFFX1 \fadd_0_0_0_0_10/n275_q_reg[7]  ( .D(\fadd_0_0_0_0_10/U29/Z_7 ), .CLK(
        clk), .QN(n13749) );
  DFFX1 \fadd_0_0_0_0_10/n280_q_reg[3]  ( .D(\fadd_0_0_0_0_10/sub_784/DIFF[3] ), .CLK(clk), .Q(\fadd_0_0_0_0_10/U4/DATA1_7 ) );
  DFFX1 \p_val_275_reg[8]  ( .D(n12430), .CLK(clk), .Q(n14038) );
  DFFX1 \p_val_297_reg[8]  ( .D(n12429), .CLK(clk), .Q(n14066) );
  DFFX1 \p_val_307_reg[8]  ( .D(n12428), .CLK(clk), .Q(n13604) );
  DFFX1 \fadd_0_0_0_0_10_x_reg[8]  ( .D(n12899), .CLK(clk), .Q(n14999), .QN(
        n12803) );
  DFFX1 \fadd_0_0_0_0_10/rightshiftercomponent/n413_q_reg[2]  ( .D(
        \fadd_0_0_0_0_10/U27/Z_2 ), .CLK(clk), .Q(
        \fadd_0_0_0_0_10/rightshiftercomponent/n44 ) );
  DFFX1 \fadd_0_0_0_0_10/rightshiftercomponent/n416_q_reg[1]  ( .D(n14973), 
        .CLK(clk), .QN(n11502) );
  DFFX1 \fadd_0_0_0_0_10/rightshiftercomponent/n416_q_reg[0]  ( .D(
        \fadd_0_0_0_0_10/rightshiftercomponent/U6/Z_0 ), .CLK(clk), .QN(n11503) );
  DFFX1 \fadd_0_0_0_0_10/rightshiftercomponent/n413_q_reg[1]  ( .D(
        \fadd_0_0_0_0_10/U27/Z_1 ), .CLK(clk), .Q(
        \fadd_0_0_0_0_10/rightshiftercomponent/n43 ) );
  DFFX1 \fadd_0_0_0_0_10/rightshiftercomponent/n417_q_reg  ( .D(
        \fadd_0_0_0_0_10/rightshiftercomponent/n11 ), .CLK(clk), .Q(n13616), 
        .QN(n11495) );
  DFFX1 \fadd_0_0_0_0_10/rightshiftercomponent/n418_q_reg[0]  ( .D(
        \fadd_0_0_0_0_10/rightshiftercomponent/U5/Z_0 ), .CLK(clk), .Q(
        \fadd_0_0_0_0_10/rightshiftercomponent/n17 ) );
  DFFX1 \fadd_0_0_0_0_10/rightshiftercomponent/n419_q_reg[0]  ( .D(
        \fadd_0_0_0_0_10/rightshiftercomponent/n17 ), .CLK(clk), .Q(
        \fadd_0_0_0_0_10/rightshiftercomponent/n16 ) );
  DFFX1 \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[5]  ( .D(
        \fadd_0_0_0_0_10/n239 ), .CLK(clk), .Q(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [5]) );
  DFFX1 \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[5]  ( .D(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [5]), .CLK(clk), 
        .Q(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/B[5] ) );
  DFFX1 \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[3]  ( .D(
        \fadd_0_0_0_0_10/n237 ), .CLK(clk), .Q(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[3]  ( .D(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [3]), .CLK(clk), 
        .Q(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/B[3] ) );
  DFFX1 \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[2]  ( .D(
        \fadd_0_0_0_0_10/n236 ), .CLK(clk), .Q(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[2]  ( .D(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [2]), .CLK(clk), 
        .Q(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/B[2] ) );
  DFFX1 \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[1]  ( .D(
        \fadd_0_0_0_0_10/n235 ), .CLK(clk), .Q(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[1]  ( .D(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [1]), .CLK(clk), 
        .Q(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/B[1] ) );
  DFFX1 \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[0]  ( .D(
        \fadd_0_0_0_0_10/n234 ), .CLK(clk), .Q(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[0]  ( .D(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [0]), .CLK(clk), 
        .Q(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/B[0] ) );
  DFFX1 \fadd_0_0_0_0_10/rightshiftercomponent/n413_q_reg[0]  ( .D(n14978), 
        .CLK(clk), .Q(\fadd_0_0_0_0_10/rightshiftercomponent/n42 ) );
  DFFX1 \fadd_0_0_0_0_10/rightshiftercomponent/n414_q_reg[0]  ( .D(
        \fadd_0_0_0_0_10/rightshiftercomponent/n42 ), .CLK(clk), .Q(
        \fadd_0_0_0_0_10/rightshiftercomponent/n41 ) );
  DFFX1 \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[4]  ( .D(
        \fadd_0_0_0_0_10/n238 ), .CLK(clk), .Q(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[4]  ( .D(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [4]), .CLK(clk), 
        .Q(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/B[4] ) );
  DFFX1 \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[6]  ( .D(
        \fadd_0_0_0_0_10/n240 ), .CLK(clk), .Q(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [6]) );
  DFFX1 \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[6]  ( .D(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [6]), .CLK(clk), 
        .Q(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/B[6] ), .QN(n13632) );
  DFFX1 \fadd_0_0_0_0_10/n278_q_reg  ( .D(n14939), .CLK(clk), .Q(
        \fadd_0_0_0_0_10/n302 ), .QN(n11497) );
  DFFX1 \fadd_0_0_0_0_10/n283_q_reg  ( .D(\fadd_0_0_0_0_10/n182 ), .CLK(clk), 
        .QN(n12069) );
  DFFX1 \p_val_275_reg[11]  ( .D(n12427), .CLK(clk), .Q(n14039) );
  DFFX1 \p_val_297_reg[11]  ( .D(n12426), .CLK(clk), .Q(n14081), .QN(n12020)
         );
  DFFX1 \p_val_307_reg[11]  ( .D(n12425), .CLK(clk), .QN(n12019) );
  DFFX1 \fadd_0_0_0_0_8_y_reg[11]  ( .D(n12884), .CLK(clk), .Q(n13501), .QN(
        n12776) );
  DFFX1 \fadd_0_0_0_0_8/n278_q_reg  ( .D(n14841), .CLK(clk), .Q(
        \fadd_0_0_0_0_8/selectclosepath_d1 ), .QN(n11594) );
  DFFX1 \fadd_0_0_0_0_8/n283_q_reg  ( .D(\fadd_0_0_0_0_8/zerofromclose ), 
        .CLK(clk), .Q(\fadd_0_0_0_0_8/zerofromclose_d1 ) );
  DFFX1 \fadd_0_0_0_0_8/n290_q_reg  ( .D(\fadd_0_0_0_0_8/ressign ), .CLK(clk), 
        .Q(\fadd_0_0_0_0_8/syncressign_d1 ) );
  DFFX1 \fadd_0_0_0_0_8/n291_q_reg  ( .D(\fadd_0_0_0_0_8/syncressign_d1 ), 
        .CLK(clk), .QN(n12017) );
  DFFX1 \p_val_227_reg[9]  ( .D(n12424), .CLK(clk), .QN(n12018) );
  DFFX1 \p_val_295_reg[9]  ( .D(n12423), .CLK(clk), .QN(n12011) );
  DFFX1 \p_val_308_reg[9]  ( .D(n12422), .CLK(clk), .QN(n12010) );
  DFFX1 \p_val_310_reg[9]  ( .D(n12421), .CLK(clk), .QN(n12008) );
  DFFX1 \fadd_0_0_0_0_8_y_reg[9]  ( .D(n12886), .CLK(clk), .QN(n11865) );
  DFFX1 \p_val_313_reg[9]  ( .D(n12420), .CLK(clk), .Q(output_p_val_313[9]) );
  DFFX1 \fadd_0_0_0_0_8_x_reg[9]  ( .D(n12874), .CLK(clk), .QN(n11877) );
  DFFX1 \fadd_0_0_0_0_8/n286_q_reg[9]  ( .D(n14848), .CLK(clk), .Q(
        \fadd_0_0_0_0_8/syncx_d1 [9]) );
  DFFX1 \fadd_0_0_0_0_8/n287_q_reg[9]  ( .D(\fadd_0_0_0_0_8/syncx_d1 [9]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_8/syncx_d2 [9]) );
  DFFX1 \fadd_0_0_0_0_8/n288_q_reg  ( .D(\fadd_0_0_0_0_8/newy_9 ), .CLK(clk), 
        .Q(\fadd_0_0_0_0_8/syncsigny_d1 ) );
  DFFX1 \fadd_0_0_0_0_8/n289_q_reg  ( .D(\fadd_0_0_0_0_8/syncsigny_d1 ), .CLK(
        clk), .QN(n12013) );
  DFFX1 \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[7]  ( .D(
        n12772), .CLK(clk), .Q(
        \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [7]) );
  DFFX1 \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[7]  ( .D(
        \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [7]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [7]) );
  DFFX1 \fadd_0_0_0_0_8/n284_q_reg  ( .D(n12772), .CLK(clk), .Q(
        \fadd_0_0_0_0_8/synceffsub_d1 ) );
  DFFX1 \fadd_0_0_0_0_8/n285_q_reg  ( .D(\fadd_0_0_0_0_8/synceffsub_d1 ), 
        .CLK(clk), .QN(n12001) );
  DFFX1 \fadd_0_0_0_0_8/n276_q_reg  ( .D(n12772), .CLK(clk), .Q(
        \fadd_0_0_0_0_8/effsub_d1 ) );
  DFFX1 \fadd_0_0_0_0_8/n277_q_reg  ( .D(\fadd_0_0_0_0_8/effsub_d1 ), .CLK(clk), .QN(n11583) );
  DFFX1 \p_val_227_reg[11]  ( .D(n12419), .CLK(clk), .QN(n12006) );
  DFFX1 \p_val_295_reg[11]  ( .D(n12418), .CLK(clk), .QN(n12005) );
  DFFX1 \p_val_308_reg[11]  ( .D(n12417), .CLK(clk), .QN(n12004) );
  DFFX1 \p_val_310_reg[11]  ( .D(n12416), .CLK(clk), .Q(n13814) );
  DFFX1 \p_val_313_reg[11]  ( .D(n12415), .CLK(clk), .Q(output_p_val_313[11])
         );
  DFFX1 \fadd_0_0_0_0_8_x_reg[11]  ( .D(n12872), .CLK(clk), .Q(n13630), .QN(
        n12774) );
  DFFX1 \fadd_0_0_0_0_8/n293_q_reg[1]  ( .D(\fadd_0_0_0_0_8/newy_11 ), .CLK(
        clk), .Q(\fadd_0_0_0_0_8/syncexnxy_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_8/n294_q_reg[1]  ( .D(\fadd_0_0_0_0_8/syncexnxy_d1 [1]), 
        .CLK(clk), .Q(n13735), .QN(n12015) );
  DFFX1 \fadd_0_0_0_0_8/n293_q_reg[3]  ( .D(\fadd_0_0_0_0_8/newx [11]), .CLK(
        clk), .Q(\fadd_0_0_0_0_8/syncexnxy_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_8/n294_q_reg[3]  ( .D(\fadd_0_0_0_0_8/syncexnxy_d1 [3]), 
        .CLK(clk), .QN(n12014) );
  DFFX1 \p_val_227_reg[10]  ( .D(n12414), .CLK(clk), .QN(n12002) );
  DFFX1 \p_val_295_reg[10]  ( .D(n12413), .CLK(clk), .QN(n12000) );
  DFFX1 \p_val_308_reg[10]  ( .D(n12412), .CLK(clk), .QN(n11999) );
  DFFX1 \p_val_310_reg[10]  ( .D(n12411), .CLK(clk), .Q(n13815) );
  DFFX1 \fadd_0_0_0_0_8_y_reg[10]  ( .D(n12885), .CLK(clk), .Q(n13588), .QN(
        n11867) );
  DFFX1 \p_val_313_reg[10]  ( .D(n12410), .CLK(clk), .Q(output_p_val_313[10])
         );
  DFFX1 \fadd_0_0_0_0_8_x_reg[10]  ( .D(n12873), .CLK(clk), .Q(n13628), .QN(
        n12775) );
  DFFX1 \fadd_0_0_0_0_8/n293_q_reg[2]  ( .D(\fadd_0_0_0_0_8/newx [10]), .CLK(
        clk), .Q(\fadd_0_0_0_0_8/syncexnxy_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_8/n294_q_reg[2]  ( .D(\fadd_0_0_0_0_8/syncexnxy_d1 [2]), 
        .CLK(clk), .Q(n13723), .QN(n12012) );
  DFFX1 \fadd_0_0_0_0_8/n293_q_reg[0]  ( .D(\fadd_0_0_0_0_8/newy_10 ), .CLK(
        clk), .Q(\fadd_0_0_0_0_8/syncexnxy_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_8/n294_q_reg[0]  ( .D(\fadd_0_0_0_0_8/syncexnxy_d1 [0]), 
        .CLK(clk), .Q(n12016) );
  DFFX1 \p_val_227_reg[2]  ( .D(n12409), .CLK(clk), .QN(n11997) );
  DFFX1 \p_val_295_reg[2]  ( .D(n12408), .CLK(clk), .QN(n11996) );
  DFFX1 \p_val_308_reg[2]  ( .D(n12407), .CLK(clk), .QN(n11995) );
  DFFX1 \p_val_310_reg[2]  ( .D(n12406), .CLK(clk), .Q(n13782) );
  DFFX1 \fadd_0_0_0_0_8_y_reg[2]  ( .D(n12893), .CLK(clk), .Q(n13593), .QN(
        n11858) );
  DFFX1 \p_val_313_reg[2]  ( .D(n12405), .CLK(clk), .Q(output_p_val_313[2]) );
  DFFX1 \fadd_0_0_0_0_8_x_reg[2]  ( .D(n12881), .CLK(clk), .QN(n11870) );
  DFFX1 \fadd_0_0_0_0_8/n286_q_reg[2]  ( .D(
        \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ), .CLK(clk), .Q(\fadd_0_0_0_0_8/syncx_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_8/n287_q_reg[2]  ( .D(\fadd_0_0_0_0_8/syncx_d1 [2]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_8/syncx_d2 [2]) );
  DFFX1 \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/n432_q_reg[4]  ( .D(
        \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ), .CLK(clk), .Q(\fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/n433_q_reg[4]  ( .D(
        \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [4]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/x_d2 [4]) );
  DFFX1 \p_val_227_reg[3]  ( .D(n12404), .CLK(clk), .QN(n11993) );
  DFFX1 \p_val_295_reg[3]  ( .D(n12403), .CLK(clk), .QN(n11992) );
  DFFX1 \p_val_308_reg[3]  ( .D(n12402), .CLK(clk), .QN(n11991) );
  DFFX1 \p_val_310_reg[3]  ( .D(n12401), .CLK(clk), .Q(n13783) );
  DFFX1 \fadd_0_0_0_0_8_y_reg[3]  ( .D(n12892), .CLK(clk), .Q(n13594), .QN(
        n11859) );
  DFFX1 \p_val_313_reg[3]  ( .D(n12400), .CLK(clk), .Q(output_p_val_313[3]) );
  DFFX1 \fadd_0_0_0_0_8_x_reg[3]  ( .D(n12880), .CLK(clk), .QN(n11871) );
  DFFX1 \fadd_0_0_0_0_8/n286_q_reg[3]  ( .D(
        \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ), .CLK(clk), .Q(\fadd_0_0_0_0_8/syncx_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_8/n287_q_reg[3]  ( .D(\fadd_0_0_0_0_8/syncx_d1 [3]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_8/syncx_d2 [3]) );
  DFFX1 \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/n432_q_reg[5]  ( .D(
        \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ), .CLK(clk), .Q(\fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [5]) );
  DFFX1 \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/n433_q_reg[5]  ( .D(
        \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [5]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/x_d2 [5]) );
  DFFX1 \p_val_227_reg[4]  ( .D(n12399), .CLK(clk), .QN(n11989) );
  DFFX1 \p_val_295_reg[4]  ( .D(n12398), .CLK(clk), .QN(n11988) );
  DFFX1 \p_val_308_reg[4]  ( .D(n12397), .CLK(clk), .QN(n11987) );
  DFFX1 \p_val_310_reg[4]  ( .D(n12396), .CLK(clk), .Q(n13784) );
  DFFX1 \fadd_0_0_0_0_8_y_reg[4]  ( .D(n12891), .CLK(clk), .Q(n5406), .QN(
        n14623) );
  DFFX1 \p_val_313_reg[4]  ( .D(n12395), .CLK(clk), .Q(output_p_val_313[4]) );
  DFFX1 \fadd_0_0_0_0_8_x_reg[4]  ( .D(n12879), .CLK(clk), .Q(n5418), .QN(
        n14628) );
  DFFX1 \fadd_0_0_0_0_8/n275_q_reg[4]  ( .D(\fadd_0_0_0_0_8/newx [4]), .CLK(
        clk), .Q(\fadd_0_0_0_0_8/newx_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_8/n281_q_reg[0]  ( .D(\fadd_0_0_0_0_8/newx [4]), .CLK(
        clk), .Q(\fadd_0_0_0_0_8/exponentresultfar0_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_8/n282_q_reg[0]  ( .D(
        \fadd_0_0_0_0_8/exponentresultfar0_d1 [0]), .CLK(clk), .Q(
        \fadd_0_0_0_0_8/exponentresultfar0_d2 [0]) );
  DFFX1 \fadd_0_0_0_0_8/n286_q_reg[4]  ( .D(\fadd_0_0_0_0_8/newx [4]), .CLK(
        clk), .Q(\fadd_0_0_0_0_8/syncx_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_8/n287_q_reg[4]  ( .D(\fadd_0_0_0_0_8/syncx_d1 [4]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_8/syncx_d2 [4]) );
  DFFX1 \p_val_227_reg[5]  ( .D(n12394), .CLK(clk), .QN(n11985) );
  DFFX1 \p_val_295_reg[5]  ( .D(n12393), .CLK(clk), .QN(n11984) );
  DFFX1 \p_val_308_reg[5]  ( .D(n12392), .CLK(clk), .QN(n11983) );
  DFFX1 \p_val_310_reg[5]  ( .D(n12391), .CLK(clk), .Q(n13785) );
  DFFX1 \fadd_0_0_0_0_8_y_reg[5]  ( .D(n12890), .CLK(clk), .Q(n5407), .QN(
        n14622) );
  DFFX1 \p_val_313_reg[5]  ( .D(n12390), .CLK(clk), .Q(output_p_val_313[5]) );
  DFFX1 \fadd_0_0_0_0_8_x_reg[5]  ( .D(n12878), .CLK(clk), .Q(n5419), .QN(
        n14627) );
  DFFX1 \fadd_0_0_0_0_8/n275_q_reg[5]  ( .D(\fadd_0_0_0_0_8/newx [5]), .CLK(
        clk), .Q(\fadd_0_0_0_0_8/newx_d1 [5]) );
  DFFX1 \fadd_0_0_0_0_8/n281_q_reg[1]  ( .D(\fadd_0_0_0_0_8/newx [5]), .CLK(
        clk), .Q(\fadd_0_0_0_0_8/exponentresultfar0_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_8/n282_q_reg[1]  ( .D(
        \fadd_0_0_0_0_8/exponentresultfar0_d1 [1]), .CLK(clk), .Q(
        \fadd_0_0_0_0_8/exponentresultfar0_d2 [1]) );
  DFFX1 \fadd_0_0_0_0_8/n286_q_reg[5]  ( .D(\fadd_0_0_0_0_8/newx [5]), .CLK(
        clk), .Q(\fadd_0_0_0_0_8/syncx_d1 [5]) );
  DFFX1 \fadd_0_0_0_0_8/n287_q_reg[5]  ( .D(\fadd_0_0_0_0_8/syncx_d1 [5]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_8/syncx_d2 [5]) );
  DFFX1 \p_val_227_reg[6]  ( .D(n12389), .CLK(clk), .QN(n11981) );
  DFFX1 \p_val_295_reg[6]  ( .D(n12388), .CLK(clk), .QN(n11980) );
  DFFX1 \p_val_308_reg[6]  ( .D(n12387), .CLK(clk), .QN(n11979) );
  DFFX1 \p_val_310_reg[6]  ( .D(n12386), .CLK(clk), .Q(n13786) );
  DFFX1 \fadd_0_0_0_0_8_y_reg[6]  ( .D(n12889), .CLK(clk), .Q(n5408), .QN(
        n14621) );
  DFFX1 \p_val_313_reg[6]  ( .D(n12385), .CLK(clk), .Q(output_p_val_313[6]) );
  DFFX1 \fadd_0_0_0_0_8_x_reg[6]  ( .D(n12877), .CLK(clk), .Q(n5420), .QN(
        n14626) );
  DFFX1 \fadd_0_0_0_0_8/n275_q_reg[6]  ( .D(\fadd_0_0_0_0_8/newx [6]), .CLK(
        clk), .Q(\fadd_0_0_0_0_8/newx_d1 [6]) );
  DFFX1 \fadd_0_0_0_0_8/n281_q_reg[2]  ( .D(\fadd_0_0_0_0_8/newx [6]), .CLK(
        clk), .Q(\fadd_0_0_0_0_8/exponentresultfar0_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_8/n282_q_reg[2]  ( .D(
        \fadd_0_0_0_0_8/exponentresultfar0_d1 [2]), .CLK(clk), .Q(
        \fadd_0_0_0_0_8/exponentresultfar0_d2 [2]) );
  DFFX1 \fadd_0_0_0_0_8/n286_q_reg[6]  ( .D(\fadd_0_0_0_0_8/newx [6]), .CLK(
        clk), .Q(\fadd_0_0_0_0_8/syncx_d1 [6]) );
  DFFX1 \fadd_0_0_0_0_8/n287_q_reg[6]  ( .D(\fadd_0_0_0_0_8/syncx_d1 [6]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_8/syncx_d2 [6]) );
  DFFX1 \p_val_227_reg[7]  ( .D(n12384), .CLK(clk), .QN(n11977) );
  DFFX1 \p_val_295_reg[7]  ( .D(n12383), .CLK(clk), .QN(n11976) );
  DFFX1 \p_val_308_reg[7]  ( .D(n12382), .CLK(clk), .QN(n11975) );
  DFFX1 \p_val_310_reg[7]  ( .D(n12381), .CLK(clk), .Q(n13787) );
  DFFX1 \fadd_0_0_0_0_8_y_reg[7]  ( .D(n12888), .CLK(clk), .Q(n5409), .QN(
        n14620) );
  DFFX1 \p_val_313_reg[7]  ( .D(n12380), .CLK(clk), .Q(output_p_val_313[7]) );
  DFFX1 \fadd_0_0_0_0_8_x_reg[7]  ( .D(n12876), .CLK(clk), .Q(n5421), .QN(
        n14625) );
  DFFX1 \fadd_0_0_0_0_8/n275_q_reg[7]  ( .D(\fadd_0_0_0_0_8/newx [7]), .CLK(
        clk), .Q(\fadd_0_0_0_0_8/newx_d1 [7]) );
  DFFX1 \fadd_0_0_0_0_8/n281_q_reg[3]  ( .D(\fadd_0_0_0_0_8/newx [7]), .CLK(
        clk), .Q(\fadd_0_0_0_0_8/exponentresultfar0_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_8/n282_q_reg[3]  ( .D(
        \fadd_0_0_0_0_8/exponentresultfar0_d1 [3]), .CLK(clk), .Q(
        \fadd_0_0_0_0_8/exponentresultfar0_d2 [3]) );
  DFFX1 \fadd_0_0_0_0_8/n286_q_reg[7]  ( .D(\fadd_0_0_0_0_8/newx [7]), .CLK(
        clk), .Q(\fadd_0_0_0_0_8/syncx_d1 [7]) );
  DFFX1 \fadd_0_0_0_0_8/n287_q_reg[7]  ( .D(\fadd_0_0_0_0_8/syncx_d1 [7]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_8/syncx_d2 [7]) );
  DFFX1 \p_val_227_reg[8]  ( .D(n12379), .CLK(clk), .QN(n11973) );
  DFFX1 \p_val_295_reg[8]  ( .D(n12378), .CLK(clk), .QN(n11972) );
  DFFX1 \p_val_308_reg[8]  ( .D(n12377), .CLK(clk), .QN(n11971) );
  DFFX1 \p_val_310_reg[8]  ( .D(n12376), .CLK(clk), .Q(n13788) );
  DFFX1 \fadd_0_0_0_0_8_y_reg[8]  ( .D(n12887), .CLK(clk), .Q(n5410), .QN(
        n14619) );
  DFFX1 \p_val_313_reg[8]  ( .D(n12375), .CLK(clk), .Q(output_p_val_313[8]) );
  DFFX1 \fadd_0_0_0_0_8_x_reg[8]  ( .D(n12875), .CLK(clk), .Q(n5422), .QN(
        n14624) );
  DFFX1 \fadd_0_0_0_0_8/rightshiftercomponent/n413_q_reg[2]  ( .D(n14842), 
        .CLK(clk), .Q(\fadd_0_0_0_0_8/rightshiftercomponent/ps_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_8/rightshiftercomponent/n416_q_reg[1]  ( .D(
        \fadd_0_0_0_0_8/rightshiftercomponent/level2[1] ), .CLK(clk), .QN(
        n11591) );
  DFFX1 \fadd_0_0_0_0_8/rightshiftercomponent/n416_q_reg[0]  ( .D(n12771), 
        .CLK(clk), .QN(n11592) );
  DFFX1 \fadd_0_0_0_0_8/rightshiftercomponent/n413_q_reg[1]  ( .D(n14845), 
        .CLK(clk), .Q(\fadd_0_0_0_0_8/rightshiftercomponent/ps_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[5]  ( .D(
        \fadd_0_0_0_0_8/fracyfarxorop [5]), .CLK(clk), .Q(
        \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [5]) );
  DFFX1 \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[5]  ( .D(
        \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [5]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [5]) );
  DFFX1 \fadd_0_0_0_0_8/rightshiftercomponent/n413_q_reg[0]  ( .D(n12769), 
        .CLK(clk), .Q(\fadd_0_0_0_0_8/rightshiftercomponent/ps_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_8/rightshiftercomponent/n414_q_reg[0]  ( .D(
        \fadd_0_0_0_0_8/rightshiftercomponent/ps_d1 [0]), .CLK(clk), .Q(
        \fadd_0_0_0_0_8/rightshiftercomponent/ps_d2[0] ) );
  DFFX1 \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[4]  ( .D(
        \fadd_0_0_0_0_8/fracyfarxorop [4]), .CLK(clk), .Q(
        \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[4]  ( .D(
        \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [4]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [4]) );
  DFFX1 \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[6]  ( .D(
        \fadd_0_0_0_0_8/fracyfarxorop [6]), .CLK(clk), .Q(
        \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [6]) );
  DFFX1 \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[6]  ( .D(
        \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [6]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [6]) );
  DFFX1 \fadd_0_0_0_0_8/n275_q_reg[8]  ( .D(\fadd_0_0_0_0_8/newx [8]), .CLK(
        clk), .Q(\fadd_0_0_0_0_8/newx_d1 [8]) );
  DFFX1 \fadd_0_0_0_0_8/n280_q_reg[0]  ( .D(
        \fadd_0_0_0_0_8/exponentresultclose [0]), .CLK(clk), .Q(
        \fadd_0_0_0_0_8/exponentresultclose_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_8/n280_q_reg[1]  ( .D(
        \fadd_0_0_0_0_8/exponentresultclose [1]), .CLK(clk), .Q(
        \fadd_0_0_0_0_8/exponentresultclose_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_8/n280_q_reg[2]  ( .D(
        \fadd_0_0_0_0_8/exponentresultclose [2]), .CLK(clk), .Q(
        \fadd_0_0_0_0_8/exponentresultclose_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_8/n280_q_reg[3]  ( .D(
        \fadd_0_0_0_0_8/exponentresultclose [3]), .CLK(clk), .Q(
        \fadd_0_0_0_0_8/exponentresultclose_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_8/n280_q_reg[4]  ( .D(
        \fadd_0_0_0_0_8/exponentresultclose [4]), .CLK(clk), .Q(
        \fadd_0_0_0_0_8/exponentresultclose_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_8/n280_q_reg[6]  ( .D(n13654), .CLK(clk), .Q(
        \fadd_0_0_0_0_8/exponentresultclose_d1 [6]) );
  DFFX1 \fadd_0_0_0_0_8/n280_q_reg[5]  ( .D(n13654), .CLK(clk), .Q(
        \fadd_0_0_0_0_8/exponentresultclose_d1 [5]) );
  DFFX1 \fadd_0_0_0_0_8/n281_q_reg[4]  ( .D(\fadd_0_0_0_0_8/newx [8]), .CLK(
        clk), .Q(\fadd_0_0_0_0_8/exponentresultfar0_d1 [4]) );
  DFFX1 \fadd_0_0_0_0_8/n282_q_reg[4]  ( .D(
        \fadd_0_0_0_0_8/exponentresultfar0_d1 [4]), .CLK(clk), .Q(
        \fadd_0_0_0_0_8/exponentresultfar0_d2 [4]) );
  DFFX1 \fadd_0_0_0_0_8/n286_q_reg[8]  ( .D(\fadd_0_0_0_0_8/newx [8]), .CLK(
        clk), .Q(\fadd_0_0_0_0_8/syncx_d1 [8]) );
  DFFX1 \fadd_0_0_0_0_8/n287_q_reg[8]  ( .D(\fadd_0_0_0_0_8/syncx_d1 [8]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_8/syncx_d2 [8]) );
  DFFX1 \p_val_227_reg[1]  ( .D(n12374), .CLK(clk), .QN(n11969) );
  DFFX1 \p_val_295_reg[1]  ( .D(n12373), .CLK(clk), .QN(n11968) );
  DFFX1 \p_val_308_reg[1]  ( .D(n12372), .CLK(clk), .QN(n11967) );
  DFFX1 \p_val_310_reg[1]  ( .D(n12371), .CLK(clk), .Q(n13789) );
  DFFX1 \fadd_0_0_0_0_8_y_reg[1]  ( .D(n12894), .CLK(clk), .Q(n13592), .QN(
        n11857) );
  DFFX1 \p_val_313_reg[1]  ( .D(n12370), .CLK(clk), .Q(output_p_val_313[1]) );
  DFFX1 \fadd_0_0_0_0_8_x_reg[1]  ( .D(n12882), .CLK(clk), .QN(n11869) );
  DFFX1 \fadd_0_0_0_0_8/rightshiftercomponent/n415_q_reg[3]  ( .D(n14851), 
        .CLK(clk), .QN(n11590) );
  DFFX1 \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[3]  ( .D(
        \fadd_0_0_0_0_8/fracyfarxorop [3]), .CLK(clk), .Q(
        \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[3]  ( .D(
        \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [3]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [3]) );
  DFFX1 \fadd_0_0_0_0_8/n286_q_reg[1]  ( .D(
        \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ), .CLK(clk), .Q(\fadd_0_0_0_0_8/syncx_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_8/n287_q_reg[1]  ( .D(\fadd_0_0_0_0_8/syncx_d1 [1]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_8/syncx_d2 [1]) );
  DFFX1 \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/n432_q_reg[3]  ( .D(
        \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ), .CLK(clk), .Q(\fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [3]) );
  DFFX1 \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/n433_q_reg[3]  ( .D(
        \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [3]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/x_d2 [3]) );
  DFFX1 \p_val_227_reg[0]  ( .D(n12369), .CLK(clk), .QN(n11965) );
  DFFX1 \p_val_295_reg[0]  ( .D(n12368), .CLK(clk), .QN(n11964) );
  DFFX1 \p_val_308_reg[0]  ( .D(n12367), .CLK(clk), .QN(n11963) );
  DFFX1 \p_val_310_reg[0]  ( .D(n12366), .CLK(clk), .Q(n13790) );
  DFFX1 \fadd_0_0_0_0_8_y_reg[0]  ( .D(n12895), .CLK(clk), .Q(n13591), .QN(
        n11856) );
  DFFX1 \p_val_313_reg[0]  ( .D(n12365), .CLK(clk), .Q(output_p_val_313[0]) );
  DFFX1 \fadd_0_0_0_0_8_x_reg[0]  ( .D(n12883), .CLK(clk), .QN(n11868) );
  DFFX1 \fadd_0_0_0_0_8/rightshiftercomponent/n415_q_reg[2]  ( .D(n14852), 
        .CLK(clk), .QN(n11589) );
  DFFX1 \fadd_0_0_0_0_8/rightshiftercomponent/n417_q_reg  ( .D(
        \fadd_0_0_0_0_8/rightshiftercomponent/n389_o ), .CLK(clk), .Q(n15002)
         );
  DFFX1 \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[2]  ( .D(
        \fadd_0_0_0_0_8/fracyfarxorop [2]), .CLK(clk), .Q(
        \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[2]  ( .D(
        \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [2]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [2]) );
  DFFX1 \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[1]  ( .D(
        \fadd_0_0_0_0_8/fracyfarxorop [1]), .CLK(clk), .Q(
        \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [1]) );
  DFFX1 \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[1]  ( .D(
        \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [1]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [1]) );
  DFFX1 \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/n434_q_reg[0]  ( .D(
        \fadd_0_0_0_0_8/fracyfarxorop [0]), .CLK(clk), .Q(
        \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/n435_q_reg[0]  ( .D(
        \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/y_d1 [0]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/y_d2 [0]) );
  DFFX1 \fadd_0_0_0_0_8/rightshiftercomponent/n418_q_reg[0]  ( .D(n12770), 
        .CLK(clk), .Q(\fadd_0_0_0_0_8/rightshiftercomponent/level1_d1[0] ) );
  DFFX1 \fadd_0_0_0_0_8/rightshiftercomponent/n419_q_reg[0]  ( .D(
        \fadd_0_0_0_0_8/rightshiftercomponent/level1_d1[0] ), .CLK(clk), .Q(
        \fadd_0_0_0_0_8/rightshiftercomponent/level1_d2[0] ) );
  DFFX1 \fadd_0_0_0_0_8/n286_q_reg[0]  ( .D(
        \add_0_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .CLK(clk), .Q(\fadd_0_0_0_0_8/syncx_d1 [0]) );
  DFFX1 \fadd_0_0_0_0_8/n287_q_reg[0]  ( .D(\fadd_0_0_0_0_8/syncx_d1 [0]), 
        .CLK(clk), .Q(\fadd_0_0_0_0_8/syncx_d2 [0]) );
  DFFX1 \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/n432_q_reg[2]  ( .D(
        \add_0_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .CLK(clk), .Q(\fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [2]) );
  DFFX1 \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/n433_q_reg[2]  ( .D(
        \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/x_d1 [2]), .CLK(clk), 
        .Q(\fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/x_d2 [2]) );
  DFFX1 \fadd_0_0_0_0_10_x_reg[11]  ( .D(n12896), .CLK(clk), .Q(n13500), .QN(
        n12802) );
  DFFX1 \fadd_0_0_0_0_10/n293_q_reg[1]  ( .D(\fadd_0_0_0_0_10/U28/Z_6 ), .CLK(
        clk), .Q(\fadd_0_0_0_0_10/n143 ) );
  DFFX1 \fadd_0_0_0_0_10/n294_q_reg[1]  ( .D(\fadd_0_0_0_0_10/n143 ), .CLK(clk), .QN(n12071) );
  DFFX1 \fadd_0_0_0_0_10/n293_q_reg[3]  ( .D(\fadd_0_0_0_0_10/U29/Z_11 ), 
        .CLK(clk), .Q(\fadd_0_0_0_0_10/n145 ) );
  DFFX1 \fadd_0_0_0_0_10/n294_q_reg[3]  ( .D(\fadd_0_0_0_0_10/n145 ), .CLK(clk), .QN(n12072) );
  DFFX1 \fadd_0_0_0_0_10/n284_q_reg  ( .D(n14938), .CLK(clk), .Q(
        \fadd_0_0_0_0_10/n169 ) );
  DFFX1 \fadd_0_0_0_0_10/n285_q_reg  ( .D(\fadd_0_0_0_0_10/n169 ), .CLK(clk), 
        .QN(n12070) );
  AO22X1 U3 ( .IN1(output_p_val_313[0]), .IN2(n12007), .IN3(n8208), .IN4(
        n13748), .Q(n12365) );
  AO22X1 U4 ( .IN1(n12009), .IN2(n13790), .IN3(n8208), .IN4(n13586), .Q(n12366) );
  OAI22X1 U6 ( .IN1(n14285), .IN2(n11964), .IN3(n14869), .IN4(n14300), .QN(
        n12368) );
  OAI22X1 U7 ( .IN1(n14266), .IN2(n11965), .IN3(n14869), .IN4(n14281), .QN(
        n12369) );
  AO22X1 U8 ( .IN1(output_p_val_313[1]), .IN2(n12007), .IN3(n8216), .IN4(
        n13748), .Q(n12370) );
  AO22X1 U9 ( .IN1(n12009), .IN2(n13789), .IN3(n8216), .IN4(n13586), .Q(n12371) );
  OAI22X1 U11 ( .IN1(n14299), .IN2(n11968), .IN3(n14868), .IN4(n14296), .QN(
        n12373) );
  OAI22X1 U12 ( .IN1(n14280), .IN2(n11969), .IN3(n14868), .IN4(n14277), .QN(
        n12374) );
  AO22X1 U13 ( .IN1(output_p_val_313[8]), .IN2(n12007), .IN3(n8219), .IN4(
        n13748), .Q(n12375) );
  AO22X1 U14 ( .IN1(n12009), .IN2(n13788), .IN3(n8219), .IN4(n13586), .Q(
        n12376) );
  OAI22X1 U16 ( .IN1(n14289), .IN2(n11972), .IN3(n14861), .IN4(n14300), .QN(
        n12378) );
  OAI22X1 U17 ( .IN1(n14270), .IN2(n11973), .IN3(n14861), .IN4(n14281), .QN(
        n12379) );
  AO22X1 U18 ( .IN1(output_p_val_313[7]), .IN2(n12007), .IN3(n8222), .IN4(
        n13748), .Q(n12380) );
  AO22X1 U19 ( .IN1(n12009), .IN2(n13787), .IN3(n8222), .IN4(n13586), .Q(
        n12381) );
  OAI22X1 U21 ( .IN1(n14217), .IN2(n11976), .IN3(n14862), .IN4(n14293), .QN(
        n12383) );
  OAI22X1 U22 ( .IN1(n14216), .IN2(n11977), .IN3(n14862), .IN4(n14274), .QN(
        n12384) );
  AO22X1 U23 ( .IN1(output_p_val_313[6]), .IN2(n12007), .IN3(n8225), .IN4(
        n13748), .Q(n12385) );
  AO22X1 U24 ( .IN1(n12009), .IN2(n13786), .IN3(n8225), .IN4(n13586), .Q(
        n12386) );
  OAI22X1 U26 ( .IN1(n14288), .IN2(n11980), .IN3(n14863), .IN4(n14223), .QN(
        n12388) );
  OAI22X1 U27 ( .IN1(n14269), .IN2(n11981), .IN3(n14863), .IN4(n14220), .QN(
        n12389) );
  AO22X1 U28 ( .IN1(output_p_val_313[5]), .IN2(n12007), .IN3(n8228), .IN4(
        n13748), .Q(n12390) );
  AO22X1 U29 ( .IN1(n12009), .IN2(n13785), .IN3(n8228), .IN4(n13586), .Q(
        n12391) );
  OAI22X1 U31 ( .IN1(n14288), .IN2(n11984), .IN3(n14864), .IN4(n14296), .QN(
        n12393) );
  OAI22X1 U32 ( .IN1(n14269), .IN2(n11985), .IN3(n14864), .IN4(n14277), .QN(
        n12394) );
  AO22X1 U33 ( .IN1(output_p_val_313[4]), .IN2(n12007), .IN3(n8231), .IN4(
        n13748), .Q(n12395) );
  AO22X1 U34 ( .IN1(n12009), .IN2(n13784), .IN3(n8231), .IN4(n13586), .Q(
        n12396) );
  OAI22X1 U36 ( .IN1(n14289), .IN2(n11988), .IN3(n14865), .IN4(n14293), .QN(
        n12398) );
  OAI22X1 U37 ( .IN1(n14270), .IN2(n11989), .IN3(n14865), .IN4(n14274), .QN(
        n12399) );
  AO22X1 U38 ( .IN1(output_p_val_313[3]), .IN2(n12007), .IN3(n8234), .IN4(
        n13748), .Q(n12400) );
  AO22X1 U39 ( .IN1(n12009), .IN2(n13783), .IN3(n8234), .IN4(n13586), .Q(
        n12401) );
  OAI22X1 U41 ( .IN1(n14290), .IN2(n11992), .IN3(n14866), .IN4(n14297), .QN(
        n12403) );
  OAI22X1 U42 ( .IN1(n14271), .IN2(n11993), .IN3(n14866), .IN4(n14278), .QN(
        n12404) );
  AO22X1 U43 ( .IN1(output_p_val_313[2]), .IN2(n12007), .IN3(n8237), .IN4(
        n13748), .Q(n12405) );
  AO22X1 U44 ( .IN1(n12009), .IN2(n13782), .IN3(n8237), .IN4(n13586), .Q(
        n12406) );
  OAI22X1 U46 ( .IN1(n14285), .IN2(n11996), .IN3(n14867), .IN4(n12356), .QN(
        n12408) );
  OAI22X1 U47 ( .IN1(n14266), .IN2(n11997), .IN3(n14867), .IN4(n12364), .QN(
        n12409) );
  AO22X1 U48 ( .IN1(output_p_val_313[10]), .IN2(n12007), .IN3(n8240), .IN4(
        n13748), .Q(n12410) );
  AO22X1 U49 ( .IN1(n12009), .IN2(n13815), .IN3(n8240), .IN4(n13586), .Q(
        n12411) );
  OAI22X1 U51 ( .IN1(n14286), .IN2(n12000), .IN3(n14860), .IN4(n14293), .QN(
        n12413) );
  OAI22X1 U52 ( .IN1(n14267), .IN2(n12002), .IN3(n14860), .IN4(n14274), .QN(
        n12414) );
  AO22X1 U53 ( .IN1(output_p_val_313[11]), .IN2(n12007), .IN3(n14858), .IN4(
        n13748), .Q(n12415) );
  AO22X1 U54 ( .IN1(n12009), .IN2(n13814), .IN3(n14858), .IN4(n13586), .Q(
        n12416) );
  OAI22X1 U57 ( .IN1(n14287), .IN2(n12005), .IN3(n8245), .IN4(n14297), .QN(
        n12418) );
  OAI22X1 U58 ( .IN1(n14268), .IN2(n12006), .IN3(n8245), .IN4(n14278), .QN(
        n12419) );
  AO22X1 U59 ( .IN1(output_p_val_313[9]), .IN2(n12007), .IN3(n15000), .IN4(
        n13748), .Q(n12420) );
  OAI22X1 U62 ( .IN1(n13586), .IN2(n12008), .IN3(n8247), .IN4(n12009), .QN(
        n12421) );
  OAI22X1 U65 ( .IN1(n14217), .IN2(n12011), .IN3(n8247), .IN4(n14294), .QN(
        n12423) );
  OAI22X1 U66 ( .IN1(n14216), .IN2(n12018), .IN3(n8247), .IN4(n14275), .QN(
        n12424) );
  OAI22X1 U67 ( .IN1(n14263), .IN2(n12019), .IN3(n12828), .IN4(n12020), .QN(
        n12425) );
  AO22X1 U68 ( .IN1(n14223), .IN2(n14081), .IN3(n8250), .IN4(n14284), .Q(
        n12426) );
  AO22X1 U70 ( .IN1(n14274), .IN2(n14039), .IN3(n8250), .IN4(n14265), .Q(
        n12427) );
  AO22X1 U71 ( .IN1(n12828), .IN2(n13604), .IN3(n14263), .IN4(n14066), .Q(
        n12428) );
  AO22X1 U72 ( .IN1(n14222), .IN2(n14066), .IN3(n8254), .IN4(n14290), .Q(
        n12429) );
  AO22X1 U74 ( .IN1(n14220), .IN2(n14038), .IN3(n8254), .IN4(n14269), .Q(
        n12430) );
  AO22X1 U75 ( .IN1(n12828), .IN2(n13603), .IN3(n14263), .IN4(n14065), .Q(
        n12431) );
  AO22X1 U76 ( .IN1(n14297), .IN2(n14065), .IN3(n8258), .IN4(n14217), .Q(
        n12432) );
  AO22X1 U78 ( .IN1(n14277), .IN2(n14037), .IN3(n8258), .IN4(n14267), .Q(
        n12433) );
  AO22X1 U79 ( .IN1(n12828), .IN2(n13602), .IN3(n14187), .IN4(n14064), .Q(
        n12434) );
  AO22X1 U80 ( .IN1(n14294), .IN2(n14064), .IN3(n8262), .IN4(n14289), .Q(
        n12435) );
  AO22X1 U82 ( .IN1(n14274), .IN2(n14036), .IN3(n8262), .IN4(n14279), .Q(
        n12436) );
  AO22X1 U83 ( .IN1(n12828), .IN2(n13601), .IN3(n14263), .IN4(n14063), .Q(
        n12437) );
  AO22X1 U84 ( .IN1(n14295), .IN2(n14063), .IN3(n8266), .IN4(n14288), .Q(
        n12438) );
  AO22X1 U86 ( .IN1(n14278), .IN2(n14035), .IN3(n8266), .IN4(n14266), .Q(
        n12439) );
  AO22X1 U87 ( .IN1(n12828), .IN2(n13600), .IN3(n14187), .IN4(n14062), .Q(
        n12440) );
  AO22X1 U88 ( .IN1(n14300), .IN2(n14062), .IN3(n8270), .IN4(n14284), .Q(
        n12441) );
  AO22X1 U90 ( .IN1(n12364), .IN2(n14034), .IN3(n8270), .IN4(n14271), .Q(
        n12442) );
  AO22X1 U91 ( .IN1(n12828), .IN2(n13599), .IN3(n14263), .IN4(n14061), .Q(
        n12443) );
  AO22X1 U92 ( .IN1(n14294), .IN2(n14061), .IN3(n8274), .IN4(n14287), .Q(
        n12444) );
  AO22X1 U134 ( .IN1(n14274), .IN2(n14033), .IN3(n8274), .IN4(n14266), .Q(
        n12445) );
  AO22X1 U135 ( .IN1(n12828), .IN2(n13598), .IN3(n14187), .IN4(n14060), .Q(
        n12446) );
  AO22X1 U136 ( .IN1(n14295), .IN2(n14060), .IN3(n8278), .IN4(n14286), .Q(
        n12447) );
  AO22X1 U138 ( .IN1(n14278), .IN2(n14032), .IN3(n8278), .IN4(n14267), .Q(
        n12448) );
  AO22X1 U139 ( .IN1(n12828), .IN2(n13597), .IN3(n14187), .IN4(n14059), .Q(
        n12449) );
  AO22X1 U140 ( .IN1(n14297), .IN2(n14059), .IN3(n8282), .IN4(n14217), .Q(
        n12450) );
  AO22X1 U142 ( .IN1(n14275), .IN2(n14031), .IN3(n8282), .IN4(n14268), .Q(
        n12451) );
  OAI22X1 U143 ( .IN1(n14187), .IN2(n12055), .IN3(n12828), .IN4(n12056), .QN(
        n12452) );
  AO22X1 U144 ( .IN1(n14295), .IN2(n14079), .IN3(n8285), .IN4(n14221), .Q(
        n12453) );
  AO22X1 U146 ( .IN1(n14277), .IN2(n14030), .IN3(n8285), .IN4(n14265), .Q(
        n12454) );
  AO22X1 U147 ( .IN1(n12828), .IN2(n13596), .IN3(n14263), .IN4(n14058), .Q(
        n12455) );
  AO22X1 U148 ( .IN1(n12356), .IN2(n14058), .IN3(n8289), .IN4(n14298), .Q(
        n12456) );
  AO22X1 U150 ( .IN1(n14219), .IN2(n14029), .IN3(n8289), .IN4(n14264), .Q(
        n12457) );
  OAI22X1 U151 ( .IN1(n14187), .IN2(n12065), .IN3(n12828), .IN4(n12066), .QN(
        n12458) );
  AO22X1 U152 ( .IN1(n14295), .IN2(n14078), .IN3(n8292), .IN4(n14285), .Q(
        n12459) );
  AO22X1 U154 ( .IN1(n14278), .IN2(n14028), .IN3(n8292), .IN4(n14270), .Q(
        n12460) );
  AO22X1 U155 ( .IN1(n14296), .IN2(n13801), .IN3(n8295), .IN4(n14290), .Q(
        n12461) );
  AO22X1 U156 ( .IN1(n14275), .IN2(n14027), .IN3(n8295), .IN4(n14271), .Q(
        n12462) );
  AO22X1 U157 ( .IN1(n14223), .IN2(n13800), .IN3(n8298), .IN4(n14301), .Q(
        n12463) );
  AO22X1 U158 ( .IN1(n14276), .IN2(n14026), .IN3(n8298), .IN4(n14266), .Q(
        n12464) );
  AO22X1 U159 ( .IN1(n14293), .IN2(n13799), .IN3(n8301), .IN4(n14217), .Q(
        n12465) );
  AO22X1 U160 ( .IN1(n14281), .IN2(n14025), .IN3(n8301), .IN4(n14216), .Q(
        n12466) );
  AO22X1 U161 ( .IN1(n14296), .IN2(n13798), .IN3(n8304), .IN4(n14283), .Q(
        n12467) );
  AO22X1 U162 ( .IN1(n14275), .IN2(n14024), .IN3(n8304), .IN4(n14273), .Q(
        n12468) );
  AO22X1 U163 ( .IN1(n14223), .IN2(n13797), .IN3(n8307), .IN4(n14285), .Q(
        n12469) );
  AO22X1 U164 ( .IN1(n14276), .IN2(n14023), .IN3(n8307), .IN4(n14264), .Q(
        n12470) );
  AO22X1 U165 ( .IN1(n14223), .IN2(n13796), .IN3(n8310), .IN4(n14290), .Q(
        n12471) );
  AO22X1 U166 ( .IN1(n14278), .IN2(n14022), .IN3(n8310), .IN4(n14270), .Q(
        n12472) );
  AO22X1 U167 ( .IN1(n14222), .IN2(n13795), .IN3(n8313), .IN4(n14289), .Q(
        n12473) );
  AO22X1 U168 ( .IN1(n14276), .IN2(n14021), .IN3(n8313), .IN4(n14268), .Q(
        n12474) );
  AO22X1 U169 ( .IN1(n14300), .IN2(n13794), .IN3(n8316), .IN4(n14288), .Q(
        n12475) );
  AO22X1 U170 ( .IN1(n12364), .IN2(n14020), .IN3(n8316), .IN4(n14218), .Q(
        n12476) );
  AO22X1 U171 ( .IN1(n14223), .IN2(n13793), .IN3(n8319), .IN4(n14284), .Q(
        n12477) );
  AO22X1 U172 ( .IN1(n14276), .IN2(n14019), .IN3(n8319), .IN4(n14267), .Q(
        n12478) );
  AO22X1 U173 ( .IN1(n14297), .IN2(n14093), .IN3(n8322), .IN4(n14292), .Q(
        n12479) );
  AO22X1 U175 ( .IN1(n14277), .IN2(n14018), .IN3(n8322), .IN4(n14216), .Q(
        n12480) );
  AO22X1 U176 ( .IN1(n14222), .IN2(n14092), .IN3(n8325), .IN4(n14291), .Q(
        n12481) );
  AO22X1 U178 ( .IN1(n14220), .IN2(n14017), .IN3(n8325), .IN4(n14282), .Q(
        n12482) );
  AO22X1 U179 ( .IN1(n14294), .IN2(n14091), .IN3(n8328), .IN4(n14287), .Q(
        n12483) );
  AO22X1 U181 ( .IN1(n14274), .IN2(n14016), .IN3(n8328), .IN4(n14280), .Q(
        n12484) );
  AO22X1 U182 ( .IN1(n12143), .IN2(n14104), .IN3(n8331), .IN4(n13587), .Q(
        n12485) );
  AO22X1 U184 ( .IN1(n14297), .IN2(n13964), .IN3(n8331), .IN4(n14288), .Q(
        n12486) );
  AO22X1 U185 ( .IN1(n14277), .IN2(n13839), .IN3(n8331), .IN4(n14282), .Q(
        n12487) );
  AO22X1 U186 ( .IN1(n12143), .IN2(n14103), .IN3(n8336), .IN4(n13587), .Q(
        n12488) );
  AO22X1 U188 ( .IN1(n14222), .IN2(n13963), .IN3(n8336), .IN4(n14301), .Q(
        n12489) );
  AO22X1 U189 ( .IN1(n14220), .IN2(n13838), .IN3(n8336), .IN4(n14280), .Q(
        n12490) );
  AO22X1 U190 ( .IN1(n12143), .IN2(n14102), .IN3(n8340), .IN4(n13587), .Q(
        n12491) );
  AO22X1 U192 ( .IN1(n12356), .IN2(n13962), .IN3(n8340), .IN4(n14217), .Q(
        n12492) );
  AO22X1 U193 ( .IN1(n14220), .IN2(n13837), .IN3(n8340), .IN4(n14216), .Q(
        n12493) );
  AO22X1 U194 ( .IN1(n12143), .IN2(n14080), .IN3(n8344), .IN4(n13587), .Q(
        n12494) );
  AO22X1 U196 ( .IN1(n14300), .IN2(n13961), .IN3(n8344), .IN4(n14298), .Q(
        n12495) );
  AO22X1 U197 ( .IN1(n14219), .IN2(n13836), .IN3(n8344), .IN4(n14282), .Q(
        n12496) );
  AO22X1 U198 ( .IN1(n12143), .IN2(n14101), .IN3(n8348), .IN4(n13587), .Q(
        n12497) );
  AO22X1 U200 ( .IN1(n14293), .IN2(n13960), .IN3(n8348), .IN4(n14283), .Q(
        n12498) );
  AO22X1 U201 ( .IN1(n14281), .IN2(n13835), .IN3(n8348), .IN4(n14267), .Q(
        n12499) );
  AO22X1 U202 ( .IN1(n12143), .IN2(n14100), .IN3(n8352), .IN4(n13587), .Q(
        n12500) );
  AO22X1 U204 ( .IN1(n14222), .IN2(n13959), .IN3(n8352), .IN4(n14284), .Q(
        n12501) );
  AO22X1 U205 ( .IN1(n14220), .IN2(n13834), .IN3(n8352), .IN4(n14216), .Q(
        n12502) );
  AO22X1 U206 ( .IN1(n12143), .IN2(n14099), .IN3(n8356), .IN4(n13587), .Q(
        n12503) );
  AO22X1 U208 ( .IN1(n14295), .IN2(n13958), .IN3(n8356), .IN4(n14292), .Q(
        n12504) );
  AO22X1 U209 ( .IN1(n14278), .IN2(n13833), .IN3(n8356), .IN4(n14271), .Q(
        n12505) );
  AO22X1 U210 ( .IN1(n12143), .IN2(n14098), .IN3(n8360), .IN4(n13587), .Q(
        n12506) );
  AO22X1 U212 ( .IN1(n12356), .IN2(n13957), .IN3(n8360), .IN4(n14291), .Q(
        n12507) );
  AO22X1 U213 ( .IN1(n14219), .IN2(n13832), .IN3(n8360), .IN4(n14282), .Q(
        n12508) );
  AO22X1 U214 ( .IN1(n12143), .IN2(n14097), .IN3(n8364), .IN4(n13587), .Q(
        n12509) );
  AO22X1 U216 ( .IN1(n14296), .IN2(n13956), .IN3(n8364), .IN4(n14217), .Q(
        n12510) );
  AO22X1 U217 ( .IN1(n14275), .IN2(n13831), .IN3(n8364), .IN4(n14270), .Q(
        n12511) );
  AO22X1 U218 ( .IN1(n12143), .IN2(n14096), .IN3(n8368), .IN4(n13587), .Q(
        n12512) );
  AO22X1 U220 ( .IN1(n14295), .IN2(n13955), .IN3(n8368), .IN4(n14292), .Q(
        n12513) );
  AO22X1 U221 ( .IN1(n14278), .IN2(n13830), .IN3(n8368), .IN4(n14265), .Q(
        n12514) );
  AO22X1 U222 ( .IN1(n12143), .IN2(n14095), .IN3(n8372), .IN4(n13587), .Q(
        n12515) );
  AO22X1 U224 ( .IN1(n12356), .IN2(n13954), .IN3(n8372), .IN4(n14291), .Q(
        n12516) );
  AO22X1 U225 ( .IN1(n14219), .IN2(n13829), .IN3(n8372), .IN4(n14264), .Q(
        n12517) );
  AO22X1 U226 ( .IN1(n12143), .IN2(n14094), .IN3(n8376), .IN4(n13587), .Q(
        n12518) );
  AO22X1 U229 ( .IN1(n14293), .IN2(n13953), .IN3(n8376), .IN4(n14217), .Q(
        n12519) );
  AO22X1 U230 ( .IN1(n12364), .IN2(n13828), .IN3(n8376), .IN4(n14216), .Q(
        n12520) );
  AO22X1 U231 ( .IN1(n14294), .IN2(n13952), .IN3(n8380), .IN4(n14221), .Q(
        n12521) );
  AO22X1 U232 ( .IN1(n14281), .IN2(n13827), .IN3(n8380), .IN4(n14282), .Q(
        n12522) );
  AO22X1 U233 ( .IN1(n14294), .IN2(n13951), .IN3(n8383), .IN4(n14298), .Q(
        n12523) );
  AO22X1 U234 ( .IN1(n14274), .IN2(n13826), .IN3(n8383), .IN4(n14280), .Q(
        n12524) );
  AO22X1 U235 ( .IN1(n12356), .IN2(n13950), .IN3(n8386), .IN4(n14299), .Q(
        n12525) );
  AO22X1 U236 ( .IN1(n14219), .IN2(n13825), .IN3(n8386), .IN4(n14279), .Q(
        n12526) );
  AO22X1 U237 ( .IN1(n14223), .IN2(n13949), .IN3(n8389), .IN4(n14283), .Q(
        n12527) );
  AO22X1 U238 ( .IN1(n14276), .IN2(n13824), .IN3(n8389), .IN4(n14279), .Q(
        n12528) );
  AO22X1 U239 ( .IN1(n14300), .IN2(n13948), .IN3(n8392), .IN4(n14292), .Q(
        n12529) );
  AO22X1 U240 ( .IN1(n12364), .IN2(n13823), .IN3(n8392), .IN4(n14218), .Q(
        n12530) );
  AO22X1 U241 ( .IN1(n14297), .IN2(n13947), .IN3(n8395), .IN4(n14217), .Q(
        n12531) );
  AO22X1 U242 ( .IN1(n14277), .IN2(n13822), .IN3(n8395), .IN4(n14272), .Q(
        n12532) );
  AO22X1 U243 ( .IN1(n14223), .IN2(n13946), .IN3(n8398), .IN4(n14221), .Q(
        n12533) );
  AO22X1 U244 ( .IN1(n14276), .IN2(n13821), .IN3(n8398), .IN4(n14280), .Q(
        n12534) );
  AO22X1 U245 ( .IN1(n14300), .IN2(n13945), .IN3(n8401), .IN4(n14299), .Q(
        n12535) );
  AO22X1 U246 ( .IN1(n12364), .IN2(n13820), .IN3(n8401), .IN4(n14279), .Q(
        n12536) );
  AO22X1 U247 ( .IN1(n14296), .IN2(n13944), .IN3(n8404), .IN4(n14287), .Q(
        n12537) );
  AO22X1 U248 ( .IN1(n14274), .IN2(n13819), .IN3(n8404), .IN4(n14268), .Q(
        n12538) );
  AO22X1 U249 ( .IN1(n14297), .IN2(n13943), .IN3(n8407), .IN4(n14286), .Q(
        n12539) );
  AO22X1 U250 ( .IN1(n14275), .IN2(n13818), .IN3(n8407), .IN4(n14273), .Q(
        n12540) );
  AO22X1 U251 ( .IN1(n14296), .IN2(n13942), .IN3(n14763), .IN4(n14221), .Q(
        n12541) );
  AO22X1 U252 ( .IN1(n14275), .IN2(n13817), .IN3(n14763), .IN4(n14266), .Q(
        n12542) );
  AO22X1 U253 ( .IN1(n14300), .IN2(n13941), .IN3(n14954), .IN4(n14298), .Q(
        n12543) );
  AO22X1 U254 ( .IN1(n12364), .IN2(n13816), .IN3(n14954), .IN4(n14280), .Q(
        n12544) );
  AO22X1 U255 ( .IN1(n14222), .IN2(n14107), .IN3(n8416), .IN4(n14299), .Q(
        n12545) );
  AO22X1 U257 ( .IN1(n14281), .IN2(n13940), .IN3(n8416), .IN4(n14271), .Q(
        n12546) );
  AO22X1 U258 ( .IN1(n14293), .IN2(n13869), .IN3(n8419), .IN4(n14301), .Q(
        n12547) );
  AO22X1 U259 ( .IN1(n14277), .IN2(n13939), .IN3(n8419), .IN4(n14218), .Q(
        n12548) );
  AO22X1 U260 ( .IN1(n14295), .IN2(n13868), .IN3(n8422), .IN4(n14217), .Q(
        n12549) );
  AO22X1 U261 ( .IN1(n14281), .IN2(n13938), .IN3(n8422), .IN4(n14272), .Q(
        n12550) );
  AO22X1 U262 ( .IN1(n14222), .IN2(n13867), .IN3(n8425), .IN4(n14283), .Q(
        n12551) );
  AO22X1 U263 ( .IN1(n14219), .IN2(n13937), .IN3(n8425), .IN4(n14216), .Q(
        n12552) );
  AO22X1 U264 ( .IN1(n14293), .IN2(n13866), .IN3(n8428), .IN4(n14284), .Q(
        n12553) );
  AO22X1 U265 ( .IN1(n14277), .IN2(n13936), .IN3(n8428), .IN4(n14273), .Q(
        n12554) );
  AO22X1 U266 ( .IN1(n14295), .IN2(n13865), .IN3(n8431), .IN4(n14287), .Q(
        n12555) );
  AO22X1 U267 ( .IN1(n14281), .IN2(n13935), .IN3(n8431), .IN4(n14269), .Q(
        n12556) );
  AO22X1 U268 ( .IN1(n14223), .IN2(n13864), .IN3(n8434), .IN4(n14286), .Q(
        n12557) );
  AO22X1 U269 ( .IN1(n14275), .IN2(n13934), .IN3(n8434), .IN4(n14270), .Q(
        n12558) );
  AO22X1 U270 ( .IN1(n14297), .IN2(n13863), .IN3(n8437), .IN4(n14284), .Q(
        n12559) );
  AO22X1 U271 ( .IN1(n14276), .IN2(n13933), .IN3(n8437), .IN4(n14216), .Q(
        n12560) );
  AO22X1 U272 ( .IN1(n14293), .IN2(n13862), .IN3(n8440), .IN4(n14291), .Q(
        n12561) );
  AO22X1 U273 ( .IN1(n12364), .IN2(n13932), .IN3(n8440), .IN4(n14273), .Q(
        n12562) );
  AO22X1 U274 ( .IN1(n12356), .IN2(n13861), .IN3(n8443), .IN4(n14283), .Q(
        n12563) );
  AO22X1 U275 ( .IN1(n14219), .IN2(n13931), .IN3(n8443), .IN4(n14269), .Q(
        n12564) );
  AO22X1 U276 ( .IN1(n14294), .IN2(n13860), .IN3(n8446), .IN4(n14298), .Q(
        n12565) );
  AO22X1 U277 ( .IN1(n14275), .IN2(n13930), .IN3(n8446), .IN4(n14218), .Q(
        n12566) );
  AO22X1 U278 ( .IN1(n14223), .IN2(n13859), .IN3(n8449), .IN4(n14301), .Q(
        n12567) );
  AO22X1 U279 ( .IN1(n12364), .IN2(n13929), .IN3(n8449), .IN4(n14272), .Q(
        n12568) );
  AO22X1 U280 ( .IN1(n14294), .IN2(n14106), .IN3(n8452), .IN4(n14217), .Q(
        n12569) );
  AO22X1 U282 ( .IN1(n14220), .IN2(n14015), .IN3(n8452), .IN4(n14282), .Q(
        n12570) );
  AO22X1 U283 ( .IN1(n14222), .IN2(n13883), .IN3(n8455), .IN4(n14221), .Q(
        n12571) );
  AO22X1 U284 ( .IN1(n14275), .IN2(n14014), .IN3(n8455), .IN4(n14279), .Q(
        n12572) );
  AO22X1 U285 ( .IN1(n12356), .IN2(n13882), .IN3(n8458), .IN4(n14288), .Q(
        n12573) );
  AO22X1 U286 ( .IN1(n12364), .IN2(n14013), .IN3(n8458), .IN4(n14264), .Q(
        n12574) );
  AO22X1 U287 ( .IN1(n14295), .IN2(n13856), .IN3(n8461), .IN4(n14292), .Q(
        n12575) );
  AO22X1 U288 ( .IN1(n14274), .IN2(n14012), .IN3(n8461), .IN4(n14216), .Q(
        n12576) );
  AO22X1 U289 ( .IN1(n14294), .IN2(n13881), .IN3(n8464), .IN4(n14291), .Q(
        n12577) );
  AO22X1 U290 ( .IN1(n14278), .IN2(n14011), .IN3(n8464), .IN4(n14265), .Q(
        n12578) );
  AO22X1 U291 ( .IN1(n14300), .IN2(n13858), .IN3(n8467), .IN4(n14289), .Q(
        n12579) );
  AO22X1 U292 ( .IN1(n14220), .IN2(n14010), .IN3(n8467), .IN4(n14267), .Q(
        n12580) );
  AO22X1 U293 ( .IN1(n14296), .IN2(n13880), .IN3(n8470), .IN4(n14288), .Q(
        n12581) );
  AO22X1 U294 ( .IN1(n14276), .IN2(n14009), .IN3(n8470), .IN4(n14268), .Q(
        n12582) );
  AO22X1 U295 ( .IN1(n14222), .IN2(n13855), .IN3(n8473), .IN4(n14292), .Q(
        n12583) );
  AO22X1 U296 ( .IN1(n14274), .IN2(n14008), .IN3(n8473), .IN4(n14265), .Q(
        n12584) );
  AO22X1 U297 ( .IN1(n14300), .IN2(n13879), .IN3(n8476), .IN4(n14291), .Q(
        n12585) );
  AO22X1 U298 ( .IN1(n14219), .IN2(n14007), .IN3(n8476), .IN4(n14264), .Q(
        n12586) );
  AO22X1 U299 ( .IN1(n14296), .IN2(n13857), .IN3(n8479), .IN4(n14217), .Q(
        n12587) );
  AO22X1 U300 ( .IN1(n14276), .IN2(n14006), .IN3(n8479), .IN4(n14216), .Q(
        n12588) );
  AO22X1 U301 ( .IN1(n14300), .IN2(n13854), .IN3(n8482), .IN4(n14221), .Q(
        n12589) );
  AO22X1 U302 ( .IN1(n14274), .IN2(n14005), .IN3(n8482), .IN4(n14282), .Q(
        n12590) );
  AO22X1 U303 ( .IN1(n14293), .IN2(n13853), .IN3(n8485), .IN4(n14290), .Q(
        n12591) );
  AO22X1 U304 ( .IN1(n14219), .IN2(n14004), .IN3(n8485), .IN4(n14280), .Q(
        n12592) );
  AO22X1 U305 ( .IN1(n12356), .IN2(n13779), .IN3(n8488), .IN4(n14299), .Q(
        n12593) );
  AO22X1 U306 ( .IN1(n14281), .IN2(n14003), .IN3(n8488), .IN4(n14279), .Q(
        n12594) );
  AO22X1 U307 ( .IN1(n14294), .IN2(n13810), .IN3(n8491), .IN4(n14285), .Q(
        n12595) );
  AO22X1 U308 ( .IN1(n14277), .IN2(n14002), .IN3(n8491), .IN4(n14218), .Q(
        n12596) );
  AO22X1 U309 ( .IN1(n14294), .IN2(n13809), .IN3(n8494), .IN4(n14292), .Q(
        n12597) );
  AO22X1 U310 ( .IN1(n14278), .IN2(n14001), .IN3(n8494), .IN4(n14267), .Q(
        n12598) );
  AO22X1 U311 ( .IN1(n14293), .IN2(n13808), .IN3(n8497), .IN4(n14287), .Q(
        n12599) );
  AO22X1 U312 ( .IN1(n14277), .IN2(n14000), .IN3(n8497), .IN4(n14268), .Q(
        n12600) );
  AO22X1 U313 ( .IN1(n12356), .IN2(n13807), .IN3(n8500), .IN4(n14298), .Q(
        n12601) );
  AO22X1 U314 ( .IN1(n14281), .IN2(n13999), .IN3(n8500), .IN4(n14280), .Q(
        n12602) );
  AO22X1 U315 ( .IN1(n14295), .IN2(n13806), .IN3(n8503), .IN4(n14299), .Q(
        n12603) );
  AO22X1 U316 ( .IN1(n14220), .IN2(n13998), .IN3(n8503), .IN4(n14218), .Q(
        n12604) );
  AO22X1 U317 ( .IN1(n14296), .IN2(n13805), .IN3(n8506), .IN4(n14217), .Q(
        n12605) );
  AO22X1 U318 ( .IN1(n14278), .IN2(n13997), .IN3(n8506), .IN4(n14216), .Q(
        n12606) );
  AO22X1 U319 ( .IN1(n12356), .IN2(n13804), .IN3(n8509), .IN4(n14221), .Q(
        n12607) );
  AO22X1 U320 ( .IN1(n14281), .IN2(n13996), .IN3(n8509), .IN4(n14273), .Q(
        n12608) );
  AO22X1 U321 ( .IN1(n14295), .IN2(n13803), .IN3(n8512), .IN4(n14298), .Q(
        n12609) );
  AO22X1 U322 ( .IN1(n14220), .IN2(n13995), .IN3(n8512), .IN4(n14264), .Q(
        n12610) );
  AO22X1 U323 ( .IN1(n14222), .IN2(n13792), .IN3(n8515), .IN4(n14298), .Q(
        n12611) );
  AO22X1 U324 ( .IN1(n12364), .IN2(n13994), .IN3(n8515), .IN4(n14280), .Q(
        n12612) );
  AO22X1 U325 ( .IN1(n14293), .IN2(n13791), .IN3(n8518), .IN4(n14299), .Q(
        n12613) );
  AO22X1 U326 ( .IN1(n14275), .IN2(n13993), .IN3(n8518), .IN4(n14279), .Q(
        n12614) );
  AO22X1 U327 ( .IN1(n14300), .IN2(n13802), .IN3(n8521), .IN4(n14301), .Q(
        n12615) );
  AO22X1 U328 ( .IN1(n14275), .IN2(n13992), .IN3(n8521), .IN4(n14218), .Q(
        n12616) );
  OAI22X1 U329 ( .IN1(n14301), .IN2(n12271), .IN3(n8523), .IN4(n14296), .QN(
        n12617) );
  AO22X1 U330 ( .IN1(n14274), .IN2(n13928), .IN3(n14944), .IN4(n14272), .Q(
        n12618) );
  AO22X1 U331 ( .IN1(n14222), .IN2(n13852), .IN3(n8527), .IN4(n14283), .Q(
        n12619) );
  AO22X1 U332 ( .IN1(n12364), .IN2(n13927), .IN3(n8527), .IN4(n14216), .Q(
        n12620) );
  AO22X1 U333 ( .IN1(n14297), .IN2(n13851), .IN3(n8530), .IN4(n14217), .Q(
        n12621) );
  AO22X1 U334 ( .IN1(n14276), .IN2(n13926), .IN3(n8530), .IN4(n14273), .Q(
        n12622) );
  AO22X1 U335 ( .IN1(n12356), .IN2(n13850), .IN3(n8533), .IN4(n14289), .Q(
        n12623) );
  AO22X1 U336 ( .IN1(n14277), .IN2(n13925), .IN3(n8533), .IN4(n14272), .Q(
        n12624) );
  AO22X1 U337 ( .IN1(n14222), .IN2(n13849), .IN3(n8536), .IN4(n14284), .Q(
        n12625) );
  AO22X1 U338 ( .IN1(n12364), .IN2(n13924), .IN3(n8536), .IN4(n14216), .Q(
        n12626) );
  AO22X1 U339 ( .IN1(n14297), .IN2(n13848), .IN3(n8539), .IN4(n14290), .Q(
        n12627) );
  AO22X1 U340 ( .IN1(n14276), .IN2(n13923), .IN3(n8539), .IN4(n14273), .Q(
        n12628) );
  AO22X1 U341 ( .IN1(n14294), .IN2(n13847), .IN3(n8542), .IN4(n14301), .Q(
        n12629) );
  AO22X1 U342 ( .IN1(n14219), .IN2(n13922), .IN3(n8542), .IN4(n14265), .Q(
        n12630) );
  AO22X1 U343 ( .IN1(n14300), .IN2(n13846), .IN3(n8545), .IN4(n14286), .Q(
        n12631) );
  AO22X1 U344 ( .IN1(n14274), .IN2(n13921), .IN3(n8545), .IN4(n14264), .Q(
        n12632) );
  AO22X1 U345 ( .IN1(n14222), .IN2(n13845), .IN3(n8548), .IN4(n14291), .Q(
        n12633) );
  AO22X1 U346 ( .IN1(n14281), .IN2(n13920), .IN3(n8548), .IN4(n14279), .Q(
        n12634) );
  AO22X1 U347 ( .IN1(n14223), .IN2(n13844), .IN3(n8551), .IN4(n14217), .Q(
        n12635) );
  AO22X1 U348 ( .IN1(n12364), .IN2(n13919), .IN3(n8551), .IN4(n14272), .Q(
        n12636) );
  AO22X1 U349 ( .IN1(n14223), .IN2(n13843), .IN3(n14710), .IN4(n14301), .Q(
        n12637) );
  AO22X1 U350 ( .IN1(n14219), .IN2(n13918), .IN3(n14710), .IN4(n14282), .Q(
        n12638) );
  AO22X1 U351 ( .IN1(n14296), .IN2(n13842), .IN3(n8557), .IN4(n14299), .Q(
        n12639) );
  AO22X1 U352 ( .IN1(n14278), .IN2(n13917), .IN3(n8557), .IN4(n14269), .Q(
        n12640) );
  AO22X1 U353 ( .IN1(n14223), .IN2(n13878), .IN3(n8560), .IN4(n14299), .Q(
        n12641) );
  AO22X1 U354 ( .IN1(n14275), .IN2(n13991), .IN3(n8560), .IN4(n14268), .Q(
        n12642) );
  AO22X1 U355 ( .IN1(n14223), .IN2(n13877), .IN3(n8563), .IN4(n14217), .Q(
        n12643) );
  AO22X1 U356 ( .IN1(n14219), .IN2(n13990), .IN3(n8563), .IN4(n14216), .Q(
        n12644) );
  AO22X1 U357 ( .IN1(n14296), .IN2(n13876), .IN3(n8566), .IN4(n14221), .Q(
        n12645) );
  AO22X1 U358 ( .IN1(n14278), .IN2(n13989), .IN3(n8566), .IN4(n14273), .Q(
        n12646) );
  AO22X1 U359 ( .IN1(n14293), .IN2(n13875), .IN3(n8569), .IN4(n14286), .Q(
        n12647) );
  AO22X1 U360 ( .IN1(n14220), .IN2(n13988), .IN3(n8569), .IN4(n14269), .Q(
        n12648) );
  AO22X1 U361 ( .IN1(n12356), .IN2(n13874), .IN3(n8572), .IN4(n14289), .Q(
        n12649) );
  AO22X1 U362 ( .IN1(n14281), .IN2(n13987), .IN3(n8572), .IN4(n14270), .Q(
        n12650) );
  AO22X1 U363 ( .IN1(n14295), .IN2(n13873), .IN3(n8575), .IN4(n14287), .Q(
        n12651) );
  AO22X1 U364 ( .IN1(n14219), .IN2(n13986), .IN3(n8575), .IN4(n14271), .Q(
        n12652) );
  AO22X1 U365 ( .IN1(n14295), .IN2(n13872), .IN3(n8578), .IN4(n14292), .Q(
        n12653) );
  AO22X1 U366 ( .IN1(n14220), .IN2(n13985), .IN3(n8578), .IN4(n14266), .Q(
        n12654) );
  AO22X1 U367 ( .IN1(n14295), .IN2(n13871), .IN3(n8581), .IN4(n14283), .Q(
        n12655) );
  AO22X1 U368 ( .IN1(n14220), .IN2(n13984), .IN3(n8581), .IN4(n14264), .Q(
        n12656) );
  AO22X1 U369 ( .IN1(n14294), .IN2(n13870), .IN3(n8584), .IN4(n14285), .Q(
        n12657) );
  AO22X1 U370 ( .IN1(n14277), .IN2(n13983), .IN3(n8584), .IN4(n14216), .Q(
        n12658) );
  AO22X1 U371 ( .IN1(n14297), .IN2(n13841), .IN3(n8587), .IN4(n14291), .Q(
        n12659) );
  AO22X1 U372 ( .IN1(n14274), .IN2(n13982), .IN3(n8587), .IN4(n14282), .Q(
        n12660) );
  AO22X1 U373 ( .IN1(n14295), .IN2(n13840), .IN3(n8590), .IN4(n14289), .Q(
        n12661) );
  AO22X1 U374 ( .IN1(n14220), .IN2(n13981), .IN3(n8590), .IN4(n14271), .Q(
        n12662) );
  AO22X1 U375 ( .IN1(n14294), .IN2(n14105), .IN3(n8593), .IN4(n14290), .Q(
        n12663) );
  AO22X1 U377 ( .IN1(n14277), .IN2(n13980), .IN3(n8593), .IN4(n14266), .Q(
        n12664) );
  AO22X1 U378 ( .IN1(n14300), .IN2(n14090), .IN3(n8596), .IN4(n14284), .Q(
        n12665) );
  AO22X1 U380 ( .IN1(n14276), .IN2(n13979), .IN3(n8596), .IN4(n14279), .Q(
        n12666) );
  AO22X1 U381 ( .IN1(n14222), .IN2(n14089), .IN3(n8599), .IN4(n14283), .Q(
        n12667) );
  AO22X1 U383 ( .IN1(n12364), .IN2(n13978), .IN3(n8599), .IN4(n14218), .Q(
        n12668) );
  AO22X1 U384 ( .IN1(n14296), .IN2(n14088), .IN3(n8602), .IN4(n14286), .Q(
        n12669) );
  AO22X1 U386 ( .IN1(n14276), .IN2(n13977), .IN3(n8602), .IN4(n14272), .Q(
        n12670) );
  AO22X1 U387 ( .IN1(n14297), .IN2(n14087), .IN3(n8605), .IN4(n14287), .Q(
        n12671) );
  AO22X1 U389 ( .IN1(n14278), .IN2(n13976), .IN3(n8605), .IN4(n14267), .Q(
        n12672) );
  AO22X1 U390 ( .IN1(n14297), .IN2(n14086), .IN3(n8608), .IN4(n14290), .Q(
        n12673) );
  AO22X1 U392 ( .IN1(n14276), .IN2(n13975), .IN3(n8608), .IN4(n14268), .Q(
        n12674) );
  AO22X1 U393 ( .IN1(n14293), .IN2(n14085), .IN3(n8611), .IN4(n14285), .Q(
        n12675) );
  AO22X1 U395 ( .IN1(n14275), .IN2(n13974), .IN3(n8611), .IN4(n14265), .Q(
        n12676) );
  AO22X1 U396 ( .IN1(n14294), .IN2(n14084), .IN3(n8614), .IN4(n14298), .Q(
        n12677) );
  AO22X1 U398 ( .IN1(n14281), .IN2(n13973), .IN3(n8614), .IN4(n14269), .Q(
        n12678) );
  AO22X1 U399 ( .IN1(n14297), .IN2(n14083), .IN3(n8617), .IN4(n14285), .Q(
        n12679) );
  AO22X1 U401 ( .IN1(n14276), .IN2(n13972), .IN3(n8617), .IN4(n14270), .Q(
        n12680) );
  AO22X1 U402 ( .IN1(n14293), .IN2(n14082), .IN3(n8620), .IN4(n14288), .Q(
        n12681) );
  AO22X1 U404 ( .IN1(n14275), .IN2(n13971), .IN3(n8620), .IN4(n14216), .Q(
        n12682) );
  AO22X1 U405 ( .IN1(n12356), .IN2(n13813), .IN3(n8623), .IN4(n14286), .Q(
        n12683) );
  AO22X1 U406 ( .IN1(n14278), .IN2(n13970), .IN3(n8623), .IN4(n14271), .Q(
        n12684) );
  AO22X1 U407 ( .IN1(n14296), .IN2(n13812), .IN3(n8626), .IN4(n14301), .Q(
        n12685) );
  AO22X1 U408 ( .IN1(n14219), .IN2(n13969), .IN3(n8626), .IN4(n14265), .Q(
        n12686) );
  AO22X1 U409 ( .IN1(n12356), .IN2(n13811), .IN3(n8629), .IN4(n14217), .Q(
        n12687) );
  AO22X1 U411 ( .IN1(n14277), .IN2(n13968), .IN3(n8629), .IN4(n14272), .Q(
        n12688) );
  NOR3X0 U423 ( .IN1(n13548), .IN2(n8632), .IN3(n8633), .QN(
        \fadd_0_0_0_0_0/sub_784/B[0] ) );
  NOR3X0 U425 ( .IN1(n13547), .IN2(n8636), .IN3(n8637), .QN(
        \fadd_0_0_0_0_1/sub_784/B[0] ) );
  NOR3X0 U427 ( .IN1(n13546), .IN2(n8640), .IN3(n8641), .QN(
        \fadd_0_0_0_0_2/sub_784/B[0] ) );
  NOR3X0 U429 ( .IN1(n13545), .IN2(n8644), .IN3(n8645), .QN(
        \fadd_0_0_0_0_3/sub_784/B[0] ) );
  NOR3X0 U431 ( .IN1(n13544), .IN2(n8648), .IN3(n8649), .QN(
        \fadd_0_0_0_0_4/sub_784/B[0] ) );
  NOR3X0 U433 ( .IN1(n13543), .IN2(n8652), .IN3(n8653), .QN(
        \fadd_0_0_0_0_5/sub_784/B[0] ) );
  NOR3X0 U435 ( .IN1(n13542), .IN2(n8656), .IN3(n8657), .QN(
        \fadd_0_0_0_0_6/sub_784/B[0] ) );
  NOR3X0 U437 ( .IN1(n13541), .IN2(n8660), .IN3(n8661), .QN(
        \fadd_0_0_0_0_7/sub_784/B[0] ) );
  NOR3X0 U439 ( .IN1(n13540), .IN2(n8664), .IN3(n8665), .QN(
        \fadd_0_0_0_0_8/sub_784/B[0] ) );
  NOR3X0 U441 ( .IN1(n13539), .IN2(n8668), .IN3(n8669), .QN(
        \fadd_0_0_0_0_9/sub_784/B[0] ) );
  OA222X1 U445 ( .IN1(n12005), .IN2(n8673), .IN3(n8245), .IN4(n8674), .IN5(
        n12004), .IN6(n14918), .Q(n8672) );
  OA21X1 U446 ( .IN1(n14123), .IN2(n14859), .IN3(n12014), .Q(n8245) );
  OA222X1 U448 ( .IN1(n11959), .IN2(n12142), .IN3(n12006), .IN4(n8679), .IN5(
        n12774), .IN6(n8680), .Q(n8671) );
  OA222X1 U450 ( .IN1(n12000), .IN2(n8673), .IN3(n14860), .IN4(n8674), .IN5(
        n11999), .IN6(n14918), .Q(n8682) );
  AO221X1 U452 ( .IN1(n8678), .IN2(n14123), .IN3(n8683), .IN4(n13723), .IN5(
        n8685), .Q(n8240) );
  NOR3X0 U455 ( .IN1(\fadd_0_0_0_0_8/resultrounded [10]), .IN2(n8683), .IN3(
        \fadd_0_0_0_0_8/zerofromclose_d1 ), .QN(n8678) );
  OA222X1 U456 ( .IN1(n11959), .IN2(n12138), .IN3(n12002), .IN4(n8679), .IN5(
        n12775), .IN6(n8680), .Q(n8681) );
  OA222X1 U458 ( .IN1(n12011), .IN2(n8673), .IN3(n8247), .IN4(n8674), .IN5(
        n12010), .IN6(n14918), .Q(n8687) );
  AO22X1 U459 ( .IN1(n12017), .IN2(n15001), .IN3(n8689), .IN4(n8683), .Q(n8247) );
  NAND4X0 U461 ( .IN1(n12012), .IN2(n12013), .IN3(n8691), .IN4(n12014), .QN(
        n8690) );
  OA222X1 U464 ( .IN1(n11959), .IN2(n12107), .IN3(n12018), .IN4(n8679), .IN5(
        n11877), .IN6(n8680), .Q(n8686) );
  OA222X1 U466 ( .IN1(n11972), .IN2(n8673), .IN3(n14861), .IN4(n8674), .IN5(
        n11971), .IN6(n14918), .Q(n8694) );
  AO22X1 U468 ( .IN1(\fadd_0_0_0_0_8/resultrounded [8]), .IN2(n15001), .IN3(
        n8683), .IN4(\fadd_0_0_0_0_8/syncx_d2 [8]), .Q(n8219) );
  OA222X1 U469 ( .IN1(n11959), .IN2(n12111), .IN3(n11973), .IN4(n8679), .IN5(
        n14624), .IN6(n8680), .Q(n8693) );
  OA222X1 U471 ( .IN1(n11976), .IN2(n8673), .IN3(n14862), .IN4(n8674), .IN5(
        n11975), .IN6(n14918), .Q(n8696) );
  AO22X1 U473 ( .IN1(\fadd_0_0_0_0_8/resultrounded [7]), .IN2(n15001), .IN3(
        n8683), .IN4(\fadd_0_0_0_0_8/syncx_d2 [7]), .Q(n8222) );
  OA222X1 U474 ( .IN1(n11959), .IN2(n12114), .IN3(n11977), .IN4(n8679), .IN5(
        n14625), .IN6(n8680), .Q(n8695) );
  OA222X1 U476 ( .IN1(n11980), .IN2(n8673), .IN3(n14863), .IN4(n8674), .IN5(
        n11979), .IN6(n14918), .Q(n8698) );
  AO22X1 U478 ( .IN1(\fadd_0_0_0_0_8/resultrounded [6]), .IN2(n15001), .IN3(
        n8683), .IN4(\fadd_0_0_0_0_8/syncx_d2 [6]), .Q(n8225) );
  OA222X1 U479 ( .IN1(n11959), .IN2(n12117), .IN3(n11981), .IN4(n8679), .IN5(
        n14626), .IN6(n8680), .Q(n8697) );
  OA222X1 U481 ( .IN1(n11984), .IN2(n8673), .IN3(n14864), .IN4(n8674), .IN5(
        n11983), .IN6(n14918), .Q(n8700) );
  AO22X1 U483 ( .IN1(\fadd_0_0_0_0_8/resultrounded [5]), .IN2(n15001), .IN3(
        n8683), .IN4(\fadd_0_0_0_0_8/syncx_d2 [5]), .Q(n8228) );
  OA222X1 U484 ( .IN1(n11959), .IN2(n12120), .IN3(n11985), .IN4(n8679), .IN5(
        n14627), .IN6(n8680), .Q(n8699) );
  OA222X1 U486 ( .IN1(n11988), .IN2(n8673), .IN3(n14865), .IN4(n8674), .IN5(
        n11987), .IN6(n14918), .Q(n8702) );
  AO22X1 U488 ( .IN1(\fadd_0_0_0_0_8/resultrounded [4]), .IN2(n15001), .IN3(
        n8683), .IN4(\fadd_0_0_0_0_8/syncx_d2 [4]), .Q(n8231) );
  OA222X1 U489 ( .IN1(n11959), .IN2(n12123), .IN3(n11989), .IN4(n8679), .IN5(
        n14628), .IN6(n8680), .Q(n8701) );
  OA222X1 U491 ( .IN1(n11992), .IN2(n8673), .IN3(n14866), .IN4(n8674), .IN5(
        n11991), .IN6(n14918), .Q(n8704) );
  AO22X1 U493 ( .IN1(\fadd_0_0_0_0_8/resultrounded [3]), .IN2(n15001), .IN3(
        n8683), .IN4(\fadd_0_0_0_0_8/syncx_d2 [3]), .Q(n8234) );
  OA222X1 U494 ( .IN1(n11959), .IN2(n12126), .IN3(n11993), .IN4(n8679), .IN5(
        n11871), .IN6(n8680), .Q(n8703) );
  OA222X1 U496 ( .IN1(n11996), .IN2(n8673), .IN3(n14867), .IN4(n8674), .IN5(
        n11995), .IN6(n14918), .Q(n8706) );
  AO22X1 U498 ( .IN1(\fadd_0_0_0_0_8/resultrounded [2]), .IN2(n15001), .IN3(
        n8683), .IN4(\fadd_0_0_0_0_8/syncx_d2 [2]), .Q(n8237) );
  OA222X1 U499 ( .IN1(n11959), .IN2(n12129), .IN3(n11997), .IN4(n8679), .IN5(
        n11870), .IN6(n8680), .Q(n8705) );
  OA222X1 U501 ( .IN1(n11968), .IN2(n8673), .IN3(n14868), .IN4(n8674), .IN5(
        n11967), .IN6(n14918), .Q(n8708) );
  AO22X1 U503 ( .IN1(\fadd_0_0_0_0_8/resultrounded [1]), .IN2(n15001), .IN3(
        n8683), .IN4(\fadd_0_0_0_0_8/syncx_d2 [1]), .Q(n8216) );
  OA222X1 U504 ( .IN1(n11959), .IN2(n12132), .IN3(n11969), .IN4(n8679), .IN5(
        n11869), .IN6(n8680), .Q(n8707) );
  OA222X1 U506 ( .IN1(n11964), .IN2(n8673), .IN3(n14869), .IN4(n8674), .IN5(
        n11963), .IN6(n14918), .Q(n8710) );
  AO22X1 U509 ( .IN1(\fadd_0_0_0_0_8/resultrounded [0]), .IN2(n15001), .IN3(
        n8683), .IN4(\fadd_0_0_0_0_8/syncx_d2 [0]), .Q(n8208) );
  OA222X1 U513 ( .IN1(n11959), .IN2(n12135), .IN3(n11965), .IN4(n8679), .IN5(
        n11868), .IN6(n8680), .Q(n8709) );
  OA222X1 U515 ( .IN1(n12097), .IN2(n8673), .IN3(n8715), .IN4(n8716), .IN5(
        n12019), .IN6(n14918), .Q(n8714) );
  NOR3X0 U517 ( .IN1(n14169), .IN2(n11960), .IN3(
        \fmul_0_0_0_0_8/expsigpostround[10] ), .QN(n8717) );
  AOI222X1 U518 ( .IN1(n13814), .IN2(n13497), .IN3(\U120/DATA1_11 ), .IN4(
        n14909), .IN5(n14906), .IN6(n13501), .QN(n8713) );
  OA222X1 U521 ( .IN1(n12094), .IN2(n8673), .IN3(n8716), .IN4(n8725), .IN5(
        n12065), .IN6(n14918), .Q(n8724) );
  AO21X1 U524 ( .IN1(n14902), .IN2(n14169), .IN3(n11961), .Q(n8726) );
  AOI222X1 U527 ( .IN1(n13815), .IN2(n13497), .IN3(\U120/DATA1_10 ), .IN4(
        n14909), .IN5(n14906), .IN6(n13588), .QN(n8723) );
  OA222X1 U530 ( .IN1(n12099), .IN2(n8673), .IN3(n11866), .IN4(n8716), .IN5(
        n12055), .IN6(n14918), .Q(n8731) );
  OA222X1 U532 ( .IN1(n12008), .IN2(n11959), .IN3(n14904), .IN4(n8679), .IN5(
        n8680), .IN6(n11865), .Q(n8730) );
  OR2X1 U534 ( .IN1(n8734), .IN2(n8735), .Q(n12887) );
  AO222X1 U535 ( .IN1(n14906), .IN2(n5410), .IN3(\U120/DATA1_8 ), .IN4(n14909), 
        .IN5(n13788), .IN6(n13497), .Q(n8735) );
  AO222X1 U538 ( .IN1(n8732), .IN2(n13604), .IN3(\U120/DATA2_8 ), .IN4(n14907), 
        .IN5(n14908), .IN6(n13801), .Q(n8734) );
  OR2X1 U541 ( .IN1(n8738), .IN2(n8739), .Q(n12888) );
  AO222X1 U542 ( .IN1(n14906), .IN2(n5409), .IN3(\U120/DATA1_7 ), .IN4(n14909), 
        .IN5(n13787), .IN6(n13497), .Q(n8739) );
  AO222X1 U545 ( .IN1(n8732), .IN2(n13603), .IN3(\U120/DATA2_7 ), .IN4(n14907), 
        .IN5(n14908), .IN6(n13800), .Q(n8738) );
  OR2X1 U548 ( .IN1(n8741), .IN2(n8742), .Q(n12889) );
  AO222X1 U549 ( .IN1(n14906), .IN2(n5408), .IN3(\U120/DATA1_6 ), .IN4(n14909), 
        .IN5(n13786), .IN6(n13497), .Q(n8742) );
  AO222X1 U552 ( .IN1(n8732), .IN2(n13602), .IN3(\U120/DATA2_6 ), .IN4(n14907), 
        .IN5(n14908), .IN6(n13799), .Q(n8741) );
  OR2X1 U555 ( .IN1(n8744), .IN2(n8745), .Q(n12890) );
  AO222X1 U556 ( .IN1(n14906), .IN2(n5407), .IN3(\U120/DATA1_5 ), .IN4(n14909), 
        .IN5(n13785), .IN6(n13497), .Q(n8745) );
  AO222X1 U559 ( .IN1(n8732), .IN2(n13601), .IN3(\U120/DATA2_5 ), .IN4(n14907), 
        .IN5(n14908), .IN6(n13798), .Q(n8744) );
  OR2X1 U562 ( .IN1(n8747), .IN2(n8748), .Q(n12891) );
  AO222X1 U563 ( .IN1(n14906), .IN2(n5406), .IN3(\U120/DATA1_4 ), .IN4(n14909), 
        .IN5(n13784), .IN6(n13497), .Q(n8748) );
  AO222X1 U566 ( .IN1(n8732), .IN2(n13600), .IN3(\U120/DATA2_4 ), .IN4(n14907), 
        .IN5(n14908), .IN6(n13797), .Q(n8747) );
  OR2X1 U569 ( .IN1(n8750), .IN2(n8751), .Q(n12892) );
  AO222X1 U570 ( .IN1(n14906), .IN2(n13594), .IN3(\U120/DATA1_3 ), .IN4(n14909), .IN5(n13783), .IN6(n13497), .Q(n8751) );
  AO222X1 U573 ( .IN1(n8732), .IN2(n13599), .IN3(\U120/DATA2_3 ), .IN4(n14907), 
        .IN5(n14908), .IN6(n13796), .Q(n8750) );
  OR2X1 U576 ( .IN1(n8753), .IN2(n8754), .Q(n12893) );
  AO222X1 U577 ( .IN1(n14906), .IN2(n13593), .IN3(\U120/DATA1_2 ), .IN4(n14909), .IN5(n13782), .IN6(n13497), .Q(n8754) );
  AO222X1 U580 ( .IN1(n8732), .IN2(n13598), .IN3(\U120/DATA2_2 ), .IN4(n14907), 
        .IN5(n14908), .IN6(n13795), .Q(n8753) );
  OR2X1 U583 ( .IN1(n8756), .IN2(n8757), .Q(n12894) );
  AO222X1 U584 ( .IN1(n14906), .IN2(n13592), .IN3(\U120/DATA1_1 ), .IN4(n14909), .IN5(n13789), .IN6(n13497), .Q(n8757) );
  AO222X1 U587 ( .IN1(n8732), .IN2(n13597), .IN3(\U120/DATA2_1 ), .IN4(n14907), 
        .IN5(n14908), .IN6(n13794), .Q(n8756) );
  OR2X1 U590 ( .IN1(n8759), .IN2(n8760), .Q(n12895) );
  AO222X1 U591 ( .IN1(n14906), .IN2(n13591), .IN3(\U120/DATA1_0 ), .IN4(n14909), .IN5(n13790), .IN6(n13497), .Q(n8760) );
  AO222X1 U597 ( .IN1(n8732), .IN2(n13596), .IN3(\U120/DATA2_0 ), .IN4(n14907), 
        .IN5(n14908), .IN6(n13793), .Q(n8759) );
  AND3X1 U603 ( .IN1(n12826), .IN2(n8680), .IN3(n11959), .Q(n8763) );
  AO222X1 U608 ( .IN1(n14433), .IN2(n13500), .IN3(n14428), .IN4(n8250), .IN5(
        n14201), .IN6(n14039), .Q(n12896) );
  OAI21X1 U610 ( .IN1(n8770), .IN2(n8771), .IN3(n12072), .QN(n8250) );
  AO222X1 U611 ( .IN1(n14213), .IN2(n13469), .IN3(n14428), .IN4(n8292), .IN5(
        n14204), .IN6(n14028), .Q(n12897) );
  AO221X1 U613 ( .IN1(n14984), .IN2(n8771), .IN3(n8774), .IN4(n13724), .IN5(
        n8776), .Q(n8292) );
  XNOR2X1 U615 ( .IN1(n8777), .IN2(n8778), .Q(n8771) );
  NAND3X0 U617 ( .IN1(n12069), .IN2(n14986), .IN3(n8780), .QN(n8770) );
  XOR2X1 U618 ( .IN1(n8781), .IN2(n8782), .Q(n8780) );
  OA22X1 U619 ( .IN1(\fadd_0_0_0_0_10/U4/DATA2_10 ), .IN2(n13527), .IN3(n12068), .IN4(\fadd_0_0_0_0_10/U4/DATA1_10 ), .Q(n8782) );
  AO221X1 U621 ( .IN1(n8784), .IN2(n14992), .IN3(n13527), .IN4(
        \fadd_0_0_0_0_10/U4/DATA1_9 ), .IN5(n14985), .Q(n8778) );
  AND3X1 U624 ( .IN1(n8789), .IN2(n8790), .IN3(n8791), .Q(n8777) );
  AO222X1 U625 ( .IN1(n14209), .IN2(n13585), .IN3(n14428), .IN4(n8285), .IN5(
        n14183), .IN6(n14030), .Q(n12898) );
  AOI22X1 U627 ( .IN1(n12057), .IN2(n14986), .IN3(n8793), .IN4(n8774), .QN(
        n8285) );
  NAND4X0 U629 ( .IN1(n12072), .IN2(n13745), .IN3(n12071), .IN4(n8796), .QN(
        n8794) );
  AO222X1 U632 ( .IN1(n14211), .IN2(n14999), .IN3(n14428), .IN4(n8254), .IN5(
        n14259), .IN6(n14038), .Q(n12899) );
  AO22X1 U634 ( .IN1(n8774), .IN2(\fadd_0_0_0_0_10/U11/DATA2_8 ), .IN3(n8798), 
        .IN4(n14986), .Q(n8254) );
  XNOR2X1 U635 ( .IN1(n8799), .IN2(n8789), .Q(n8798) );
  NAND3X0 U636 ( .IN1(n8800), .IN2(n8787), .IN3(n8801), .QN(n8789) );
  OA22X1 U637 ( .IN1(n12067), .IN2(n8802), .IN3(n12024), .IN4(n12068), .Q(
        n8801) );
  OA22X1 U638 ( .IN1(n8803), .IN2(n8804), .IN3(n14987), .IN4(n8805), .Q(n8802)
         );
  NAND3X0 U639 ( .IN1(n14987), .IN2(n14994), .IN3(n12067), .QN(n8787) );
  NAND3X0 U640 ( .IN1(n14992), .IN2(n8804), .IN3(n12067), .QN(n8800) );
  AO222X1 U642 ( .IN1(n14211), .IN2(n14998), .IN3(n14428), .IN4(n8258), .IN5(
        n14183), .IN6(n14037), .Q(n12900) );
  AO22X1 U644 ( .IN1(n8774), .IN2(\fadd_0_0_0_0_10/U11/DATA2_7 ), .IN3(n8808), 
        .IN4(n14986), .Q(n8258) );
  XOR2X1 U645 ( .IN1(n8790), .IN2(n8791), .Q(n8808) );
  AO221X1 U647 ( .IN1(n8811), .IN2(n12068), .IN3(n8812), .IN4(n13722), .IN5(
        n8814), .Q(n8790) );
  AO22X1 U648 ( .IN1(n13527), .IN2(\fadd_0_0_0_0_10/U4/DATA1_7 ), .IN3(n8815), 
        .IN4(n12028), .Q(n8814) );
  AO21X1 U650 ( .IN1(n14994), .IN2(n14988), .IN3(n8817), .Q(n8812) );
  OA21X1 U652 ( .IN1(n12028), .IN2(n14988), .IN3(n8819), .Q(n8818) );
  NAND3X0 U653 ( .IN1(n14988), .IN2(n14993), .IN3(n12028), .QN(n8819) );
  AO222X1 U654 ( .IN1(n14211), .IN2(n14997), .IN3(n14428), .IN4(n8262), .IN5(
        n14916), .IN6(n14036), .Q(n12901) );
  AO22X1 U656 ( .IN1(n8774), .IN2(\fadd_0_0_0_0_10/U11/DATA2_6 ), .IN3(n8822), 
        .IN4(n14986), .Q(n8262) );
  XOR2X1 U657 ( .IN1(n8809), .IN2(n8810), .Q(n8822) );
  AOI221X1 U658 ( .IN1(n8817), .IN2(n14988), .IN3(n13527), .IN4(
        \fadd_0_0_0_0_10/U4/DATA1_6 ), .IN5(n8823), .QN(n8810) );
  AO21X1 U659 ( .IN1(n8824), .IN2(n13706), .IN3(n8815), .Q(n8823) );
  NOR3X0 U660 ( .IN1(n8805), .IN2(n14988), .IN3(n13706), .QN(n8815) );
  AO22X1 U661 ( .IN1(n14994), .IN2(n14988), .IN3(n14992), .IN4(n8826), .Q(
        n8824) );
  AO222X1 U666 ( .IN1(n14210), .IN2(n14996), .IN3(n14428), .IN4(n8266), .IN5(
        n14916), .IN6(n14035), .Q(n12902) );
  AO22X1 U668 ( .IN1(n8774), .IN2(\fadd_0_0_0_0_10/U11/DATA2_5 ), .IN3(n8830), 
        .IN4(n14986), .Q(n8266) );
  XOR2X1 U669 ( .IN1(n8828), .IN2(n8827), .Q(n8830) );
  OAI221X1 U671 ( .IN1(n8803), .IN2(n8833), .IN3(n8834), .IN4(n13677), .IN5(
        n8836), .QN(n8828) );
  OA22X1 U672 ( .IN1(n8805), .IN2(n8837), .IN3(n12037), .IN4(n12068), .Q(n8836) );
  OA22X1 U673 ( .IN1(n12041), .IN2(n8838), .IN3(n8839), .IN4(n8805), .Q(n8834)
         );
  OR2X1 U674 ( .IN1(n8839), .IN2(n12036), .Q(n8833) );
  AO222X1 U676 ( .IN1(n14208), .IN2(n13635), .IN3(n14428), .IN4(n8270), .IN5(
        n14262), .IN6(n14034), .Q(n12903) );
  OAI22X1 U678 ( .IN1(n12042), .IN2(n14986), .IN3(n8841), .IN4(n8774), .QN(
        n8270) );
  OA222X1 U679 ( .IN1(n14991), .IN2(n8842), .IN3(n14991), .IN4(n8843), .IN5(
        n8831), .IN6(n8844), .Q(n8841) );
  NAND3X0 U680 ( .IN1(n8845), .IN2(n8846), .IN3(n8842), .QN(n8831) );
  AND2X1 U681 ( .IN1(n8845), .IN2(n8846), .Q(n8843) );
  AO222X1 U683 ( .IN1(n8847), .IN2(n13697), .IN3(n8849), .IN4(n12041), .IN5(
        n13527), .IN6(\fadd_0_0_0_0_10/U4/DATA1_4 ), .Q(n8844) );
  AO222X1 U686 ( .IN1(n14212), .IN2(n13562), .IN3(n14428), .IN4(n8274), .IN5(
        n14261), .IN6(n14033), .Q(n12904) );
  AO22X1 U688 ( .IN1(n8774), .IN2(\fadd_0_0_0_0_10/U11/DATA2_3 ), .IN3(n8852), 
        .IN4(n14986), .Q(n8274) );
  XNOR2X1 U689 ( .IN1(n8853), .IN2(n8845), .Q(n8852) );
  AO221X1 U690 ( .IN1(n8847), .IN2(\fadd_0_0_0_0_10/U21/DATA2_2 ), .IN3(
        \fadd_0_0_0_0_10/U22/DATA1_3 ), .IN4(n14994), .IN5(n8854), .Q(n8845)
         );
  AO222X1 U691 ( .IN1(n8855), .IN2(\fadd_0_0_0_0_10/norm/U4/DATA2_5 ), .IN3(
        n8856), .IN4(n13695), .IN5(n14990), .IN6(\fadd_0_0_0_0_10/U21/DATA2_3 ), .Q(n8854) );
  AO222X1 U693 ( .IN1(n14433), .IN2(n13538), .IN3(n14428), .IN4(n8278), .IN5(
        n14260), .IN6(n14032), .Q(n12905) );
  AO22X1 U695 ( .IN1(n8774), .IN2(\fadd_0_0_0_0_10/U11/DATA2_2 ), .IN3(n8860), 
        .IN4(n14986), .Q(n8278) );
  XOR2X1 U696 ( .IN1(n8846), .IN2(n8842), .Q(n8860) );
  AO221X1 U698 ( .IN1(\fadd_0_0_0_0_10/U22/DATA1_3 ), .IN2(n8847), .IN3(
        \fadd_0_0_0_0_10/U22/DATA1_2 ), .IN4(n14994), .IN5(n8863), .Q(n8846)
         );
  AO222X1 U699 ( .IN1(n8855), .IN2(n13695), .IN3(n8856), .IN4(n13549), .IN5(
        \fadd_0_0_0_0_10/U21/DATA2_2 ), .IN6(n14990), .Q(n8863) );
  AO222X1 U701 ( .IN1(n14211), .IN2(n13526), .IN3(n14428), .IN4(n8282), .IN5(
        n14202), .IN6(n14031), .Q(n12906) );
  AO22X1 U703 ( .IN1(n8774), .IN2(\fadd_0_0_0_0_10/U11/DATA2_1 ), .IN3(n8866), 
        .IN4(n14986), .Q(n8282) );
  XOR2X1 U704 ( .IN1(n8861), .IN2(n8862), .Q(n8866) );
  AOI221X1 U705 ( .IN1(\fadd_0_0_0_0_10/U22/DATA1_2 ), .IN2(n8847), .IN3(
        \fadd_0_0_0_0_10/U22/DATA1_1 ), .IN4(n14994), .IN5(n8867), .QN(n8862)
         );
  AO222X1 U706 ( .IN1(n8855), .IN2(n13549), .IN3(n8856), .IN4(n13485), .IN5(
        \fadd_0_0_0_0_10/U22/DATA1_3 ), .IN6(n14990), .Q(n8867) );
  AND2X1 U710 ( .IN1(n8850), .IN2(n12068), .Q(n8847) );
  AO222X1 U712 ( .IN1(n14214), .IN2(n13477), .IN3(n14428), .IN4(n8289), .IN5(
        n14259), .IN6(n14029), .Q(n12907) );
  AO22X1 U714 ( .IN1(n8774), .IN2(\fadd_0_0_0_0_10/U11/DATA2_0 ), .IN3(n14986), 
        .IN4(n8873), .Q(n8289) );
  XOR2X1 U715 ( .IN1(n8870), .IN2(n8871), .Q(n8873) );
  AO221X1 U716 ( .IN1(n12068), .IN2(n8874), .IN3(\fadd_0_0_0_0_10/U22/DATA1_0 ), .IN4(n14994), .IN5(n8875), .Q(n8871) );
  AO22X1 U717 ( .IN1(n8855), .IN2(n13485), .IN3(n8856), .IN4(n13676), .Q(n8875) );
  AO22X1 U721 ( .IN1(n8877), .IN2(n8878), .IN3(n8879), .IN4(n8855), .Q(n8870)
         );
  AND2X1 U722 ( .IN1(n12061), .IN2(n13527), .Q(n8855) );
  NAND3X0 U725 ( .IN1(n11495), .IN2(n14989), .IN3(n8881), .QN(n8878) );
  AOI221X1 U726 ( .IN1(n14993), .IN2(\fadd_0_0_0_0_10/U20/DATA1_0 ), .IN3(
        n8882), .IN4(\fadd_0_0_0_0_10/U22/DATA1_0 ), .IN5(n8883), .QN(n8881)
         );
  OR2X1 U727 ( .IN1(n8869), .IN2(n13412), .Q(n8882) );
  AO22X1 U729 ( .IN1(\fadd_0_0_0_0_10/U22/DATA1_1 ), .IN2(n8850), .IN3(
        \fadd_0_0_0_0_10/U22/DATA1_2 ), .IN4(n8869), .Q(n8874) );
  AO22X1 U730 ( .IN1(\fadd_0_0_0_0_10/U20/DATA1_0 ), .IN2(n14994), .IN3(n12068), .IN4(n8884), .Q(n8877) );
  AO22X1 U731 ( .IN1(\fadd_0_0_0_0_10/U22/DATA1_0 ), .IN2(n8850), .IN3(
        \fadd_0_0_0_0_10/U22/DATA1_1 ), .IN4(n8869), .Q(n8884) );
  NAND4X0 U736 ( .IN1(n12071), .IN2(n12072), .IN3(n12073), .IN4(n13724), .QN(
        n8774) );
  AO222X1 U738 ( .IN1(n14209), .IN2(n13886), .IN3(n14422), .IN4(n8887), .IN5(
        \U5/DATA1_11 ), .IN6(n14262), .Q(n12908) );
  AO222X1 U743 ( .IN1(n14434), .IN2(n13887), .IN3(n8893), .IN4(n14423), .IN5(
        \U5/DATA1_10 ), .IN6(n14183), .Q(n12909) );
  OA21X1 U744 ( .IN1(n8894), .IN2(n11958), .IN3(n13771), .Q(n8893) );
  AO222X1 U747 ( .IN1(n14207), .IN2(n13726), .IN3(n14422), .IN4(\U5/DATA2_9 ), 
        .IN5(\U5/DATA1_9 ), .IN6(n14916), .Q(n12910) );
  AO222X1 U748 ( .IN1(n14433), .IN2(n14983), .IN3(n13444), .IN4(n14423), .IN5(
        p___constant_11xf32_10[8]), .IN6(n14259), .Q(n12911) );
  AO222X1 U749 ( .IN1(n14209), .IN2(n14982), .IN3(n13445), .IN4(n14423), .IN5(
        p___constant_11xf32_10[7]), .IN6(n14206), .Q(n12912) );
  AO222X1 U750 ( .IN1(n14434), .IN2(n14981), .IN3(n13446), .IN4(n14423), .IN5(
        p___constant_11xf32_10[6]), .IN6(n14201), .Q(n12913) );
  AO222X1 U751 ( .IN1(n14433), .IN2(n14980), .IN3(n13447), .IN4(n14423), .IN5(
        p___constant_11xf32_10[5]), .IN6(n14260), .Q(n12914) );
  AO222X1 U752 ( .IN1(n14214), .IN2(n13885), .IN3(n13448), .IN4(n14423), .IN5(
        p___constant_11xf32_10[4]), .IN6(n14203), .Q(n12915) );
  AO222X1 U753 ( .IN1(n14434), .IN2(n13696), .IN3(n13449), .IN4(n14423), .IN5(
        p___constant_11xf32_10[3]), .IN6(n14259), .Q(n12916) );
  AO222X1 U754 ( .IN1(n14209), .IN2(n13673), .IN3(n13450), .IN4(n14424), .IN5(
        p___constant_11xf32_10[2]), .IN6(n14201), .Q(n12917) );
  AO222X1 U755 ( .IN1(n8766), .IN2(n13646), .IN3(n13451), .IN4(n14423), .IN5(
        p___constant_11xf32_10[1]), .IN6(n14205), .Q(n12918) );
  AO222X1 U756 ( .IN1(n14207), .IN2(n13633), .IN3(n13452), .IN4(n14423), .IN5(
        p___constant_11xf32_10[0]), .IN6(n14205), .Q(n12919) );
  AO222X1 U757 ( .IN1(n14212), .IN2(n13513), .IN3(n14429), .IN4(n8325), .IN5(
        n14201), .IN6(n14017), .Q(n12920) );
  AO21X1 U759 ( .IN1(\fadd_0_0_0_0_9/resultrounded [9]), .IN2(n8906), .IN3(
        n13776), .Q(n8325) );
  AO222X1 U761 ( .IN1(n14212), .IN2(n13504), .IN3(n14429), .IN4(n8322), .IN5(
        n14262), .IN6(n14018), .Q(n12921) );
  AO221X1 U763 ( .IN1(n8906), .IN2(n14890), .IN3(n8910), .IN4(n13732), .IN5(
        n8912), .Q(n8322) );
  NOR3X0 U766 ( .IN1(\fadd_0_0_0_0_9/resultrounded [10]), .IN2(n8910), .IN3(
        \fadd_0_0_0_0_9/zerofromclose_d1 ), .QN(n8906) );
  AO222X1 U767 ( .IN1(n14207), .IN2(n13583), .IN3(n14429), .IN4(n8328), .IN5(
        n14204), .IN6(n14016), .Q(n12922) );
  AOI22X1 U769 ( .IN1(n12105), .IN2(n14959), .IN3(n8915), .IN4(n8910), .QN(
        n8328) );
  NAND4X0 U771 ( .IN1(n12100), .IN2(n12101), .IN3(n8917), .IN4(n12102), .QN(
        n8916) );
  AO222X1 U774 ( .IN1(n8766), .IN2(n5350), .IN3(n14429), .IN4(n8295), .IN5(
        n14916), .IN6(n14027), .Q(n12923) );
  AO22X1 U776 ( .IN1(\fadd_0_0_0_0_9/resultrounded [8]), .IN2(n14959), .IN3(
        n8910), .IN4(\fadd_0_0_0_0_9/syncx_d2 [8]), .Q(n8295) );
  AO222X1 U777 ( .IN1(n14210), .IN2(n5349), .IN3(n14429), .IN4(n8298), .IN5(
        n14262), .IN6(n14026), .Q(n12924) );
  AO22X1 U779 ( .IN1(\fadd_0_0_0_0_9/resultrounded [7]), .IN2(n14959), .IN3(
        n8910), .IN4(\fadd_0_0_0_0_9/syncx_d2 [7]), .Q(n8298) );
  AO222X1 U780 ( .IN1(n14209), .IN2(n5348), .IN3(n14429), .IN4(n8301), .IN5(
        n14261), .IN6(n14025), .Q(n12925) );
  AO22X1 U782 ( .IN1(\fadd_0_0_0_0_9/resultrounded [6]), .IN2(n14959), .IN3(
        n8910), .IN4(\fadd_0_0_0_0_9/syncx_d2 [6]), .Q(n8301) );
  AO222X1 U783 ( .IN1(n14213), .IN2(n5347), .IN3(n14429), .IN4(n8304), .IN5(
        n14260), .IN6(n14024), .Q(n12926) );
  AO22X1 U785 ( .IN1(\fadd_0_0_0_0_9/resultrounded [5]), .IN2(n14959), .IN3(
        n8910), .IN4(\fadd_0_0_0_0_9/syncx_d2 [5]), .Q(n8304) );
  AO222X1 U786 ( .IN1(n14433), .IN2(n5346), .IN3(n14429), .IN4(n8307), .IN5(
        n14201), .IN6(n14023), .Q(n12927) );
  AO22X1 U788 ( .IN1(\fadd_0_0_0_0_9/resultrounded [4]), .IN2(n14959), .IN3(
        n8910), .IN4(\fadd_0_0_0_0_9/syncx_d2 [4]), .Q(n8307) );
  AO222X1 U789 ( .IN1(n14212), .IN2(n13574), .IN3(n14429), .IN4(n8310), .IN5(
        n14262), .IN6(n14022), .Q(n12928) );
  AO22X1 U791 ( .IN1(\fadd_0_0_0_0_9/resultrounded [3]), .IN2(n14959), .IN3(
        n8910), .IN4(\fadd_0_0_0_0_9/syncx_d2 [3]), .Q(n8310) );
  AO222X1 U792 ( .IN1(n14214), .IN2(n13557), .IN3(n14429), .IN4(n8313), .IN5(
        n14262), .IN6(n14021), .Q(n12929) );
  AO22X1 U794 ( .IN1(\fadd_0_0_0_0_9/resultrounded [2]), .IN2(n14959), .IN3(
        n8910), .IN4(\fadd_0_0_0_0_9/syncx_d2 [2]), .Q(n8313) );
  AO222X1 U795 ( .IN1(n14208), .IN2(n13532), .IN3(n14429), .IN4(n8316), .IN5(
        n14206), .IN6(n14020), .Q(n12930) );
  AO22X1 U797 ( .IN1(\fadd_0_0_0_0_9/resultrounded [1]), .IN2(n14959), .IN3(
        n8910), .IN4(\fadd_0_0_0_0_9/syncx_d2 [1]), .Q(n8316) );
  AO222X1 U798 ( .IN1(n14214), .IN2(n13521), .IN3(n14429), .IN4(n8319), .IN5(
        n14261), .IN6(n14019), .Q(n12931) );
  AO22X1 U800 ( .IN1(\fadd_0_0_0_0_9/resultrounded [0]), .IN2(n14959), .IN3(
        n8910), .IN4(\fadd_0_0_0_0_9/syncx_d2 [0]), .Q(n8319) );
  AO222X1 U804 ( .IN1(n14213), .IN2(n13626), .IN3(n14422), .IN4(n8929), .IN5(
        \U58/DATA1_11 ), .IN6(n14183), .Q(n12932) );
  AO222X1 U809 ( .IN1(n14214), .IN2(n13893), .IN3(n8935), .IN4(n14423), .IN5(
        \U58/DATA1_10 ), .IN6(n14202), .Q(n12933) );
  OA21X1 U810 ( .IN1(n8936), .IN2(n11956), .IN3(n13770), .Q(n8935) );
  AO222X1 U813 ( .IN1(n14209), .IN2(n13721), .IN3(n14422), .IN4(\U58/DATA2_9 ), 
        .IN5(\U58/DATA1_9 ), .IN6(n14204), .Q(n12934) );
  AO222X1 U814 ( .IN1(n14210), .IN2(n5338), .IN3(\U58/DATA2_8 ), .IN4(n14424), 
        .IN5(\U58/DATA1_8 ), .IN6(n14916), .Q(n12935) );
  AO222X1 U815 ( .IN1(n14213), .IN2(n5337), .IN3(\U58/DATA2_7 ), .IN4(n14423), 
        .IN5(\U58/DATA1_7 ), .IN6(n14183), .Q(n12936) );
  AO222X1 U816 ( .IN1(n14211), .IN2(n5336), .IN3(\U58/DATA2_6 ), .IN4(n14423), 
        .IN5(\U58/DATA1_6 ), .IN6(n14203), .Q(n12937) );
  AO222X1 U817 ( .IN1(n14210), .IN2(n5335), .IN3(\U58/DATA2_5 ), .IN4(n14425), 
        .IN5(\U58/DATA1_5 ), .IN6(n14261), .Q(n12938) );
  AO222X1 U818 ( .IN1(n14208), .IN2(n5334), .IN3(\U58/DATA2_4 ), .IN4(n14424), 
        .IN5(\U58/DATA1_4 ), .IN6(n14202), .Q(n12939) );
  AO222X1 U819 ( .IN1(n14208), .IN2(n13712), .IN3(n13453), .IN4(n14424), .IN5(
        p___constant_11xf32_9[3]), .IN6(n14203), .Q(n12940) );
  AO222X1 U820 ( .IN1(n14208), .IN2(n13690), .IN3(n13454), .IN4(n14424), .IN5(
        p___constant_11xf32_9[2]), .IN6(n14260), .Q(n12941) );
  AO222X1 U821 ( .IN1(n14212), .IN2(n13669), .IN3(n13455), .IN4(n14424), .IN5(
        p___constant_11xf32_9[1]), .IN6(n14203), .Q(n12942) );
  AO222X1 U822 ( .IN1(n14208), .IN2(n13641), .IN3(n13456), .IN4(n14424), .IN5(
        p___constant_11xf32_9[0]), .IN6(n14206), .Q(n12943) );
  AO221X1 U823 ( .IN1(n8947), .IN2(n8376), .IN3(n14911), .IN4(n13953), .IN5(
        n8949), .Q(n12944) );
  AO22X1 U824 ( .IN1(n14910), .IN2(n13515), .IN3(n14420), .IN4(n13828), .Q(
        n8949) );
  AO21X1 U827 ( .IN1(\fadd_0_0_0_0_0/resultrounded [9]), .IN2(n8953), .IN3(
        n13778), .Q(n8376) );
  AO221X1 U829 ( .IN1(n8947), .IN2(n8372), .IN3(n14911), .IN4(n13954), .IN5(
        n8955), .Q(n12945) );
  AO22X1 U830 ( .IN1(n14910), .IN2(n13506), .IN3(n14420), .IN4(n13829), .Q(
        n8955) );
  AO221X1 U833 ( .IN1(n8953), .IN2(n14668), .IN3(n8958), .IN4(n13729), .IN5(
        n8960), .Q(n8372) );
  NOR3X0 U836 ( .IN1(\fadd_0_0_0_0_0/resultrounded [10]), .IN2(n8958), .IN3(
        \fadd_0_0_0_0_0/zerofromclose_d1 ), .QN(n8953) );
  AO221X1 U837 ( .IN1(n8331), .IN2(n8947), .IN3(n14911), .IN4(n13964), .IN5(
        n8961), .Q(n12946) );
  AO22X1 U838 ( .IN1(n14910), .IN2(n13595), .IN3(n14421), .IN4(n13839), .Q(
        n8961) );
  AOI22X1 U842 ( .IN1(n12109), .IN2(n14957), .IN3(n8964), .IN4(n8958), .QN(
        n8331) );
  NAND4X0 U844 ( .IN1(n12148), .IN2(n13742), .IN3(n12146), .IN4(n8967), .QN(
        n8965) );
  AO221X1 U847 ( .IN1(n8947), .IN2(n8336), .IN3(n14911), .IN4(n13963), .IN5(
        n8968), .Q(n12947) );
  AO22X1 U848 ( .IN1(n14910), .IN2(n5998), .IN3(n14421), .IN4(n13838), .Q(
        n8968) );
  AO22X1 U851 ( .IN1(\fadd_0_0_0_0_0/resultrounded [8]), .IN2(n14957), .IN3(
        n8958), .IN4(\fadd_0_0_0_0_0/syncx_d2 [8]), .Q(n8336) );
  AO221X1 U852 ( .IN1(n8947), .IN2(n8340), .IN3(n14911), .IN4(n13962), .IN5(
        n8970), .Q(n12948) );
  AO22X1 U853 ( .IN1(n14910), .IN2(n5997), .IN3(n14421), .IN4(n13837), .Q(
        n8970) );
  AO22X1 U856 ( .IN1(\fadd_0_0_0_0_0/resultrounded [7]), .IN2(n14957), .IN3(
        n8958), .IN4(\fadd_0_0_0_0_0/syncx_d2 [7]), .Q(n8340) );
  AO221X1 U857 ( .IN1(n8947), .IN2(n8344), .IN3(n14911), .IN4(n13961), .IN5(
        n8972), .Q(n12949) );
  AO22X1 U858 ( .IN1(n14910), .IN2(n5996), .IN3(n14421), .IN4(n13836), .Q(
        n8972) );
  AO22X1 U861 ( .IN1(\fadd_0_0_0_0_0/resultrounded [6]), .IN2(n14957), .IN3(
        n8958), .IN4(\fadd_0_0_0_0_0/syncx_d2 [6]), .Q(n8344) );
  AO221X1 U862 ( .IN1(n8947), .IN2(n8348), .IN3(n14911), .IN4(n13960), .IN5(
        n8974), .Q(n12950) );
  AO22X1 U863 ( .IN1(n14910), .IN2(n5995), .IN3(n14421), .IN4(n13835), .Q(
        n8974) );
  AO22X1 U866 ( .IN1(\fadd_0_0_0_0_0/resultrounded [5]), .IN2(n14957), .IN3(
        n8958), .IN4(\fadd_0_0_0_0_0/syncx_d2 [5]), .Q(n8348) );
  AO221X1 U867 ( .IN1(n8947), .IN2(n8352), .IN3(n14911), .IN4(n13959), .IN5(
        n8976), .Q(n12951) );
  AO22X1 U868 ( .IN1(n14910), .IN2(n5994), .IN3(n14420), .IN4(n13834), .Q(
        n8976) );
  AO22X1 U871 ( .IN1(\fadd_0_0_0_0_0/resultrounded [4]), .IN2(n14957), .IN3(
        n8958), .IN4(\fadd_0_0_0_0_0/syncx_d2 [4]), .Q(n8352) );
  AO221X1 U872 ( .IN1(n8947), .IN2(n8356), .IN3(n14911), .IN4(n13958), .IN5(
        n8978), .Q(n12952) );
  AO22X1 U873 ( .IN1(n14910), .IN2(n13576), .IN3(n14421), .IN4(n13833), .Q(
        n8978) );
  AO22X1 U876 ( .IN1(\fadd_0_0_0_0_0/resultrounded [3]), .IN2(n14957), .IN3(
        n8958), .IN4(\fadd_0_0_0_0_0/syncx_d2 [3]), .Q(n8356) );
  AO221X1 U877 ( .IN1(n8947), .IN2(n8360), .IN3(n14911), .IN4(n13957), .IN5(
        n8980), .Q(n12953) );
  AO22X1 U878 ( .IN1(n14910), .IN2(n13559), .IN3(n14421), .IN4(n13832), .Q(
        n8980) );
  AO22X1 U881 ( .IN1(\fadd_0_0_0_0_0/resultrounded [2]), .IN2(n14957), .IN3(
        n8958), .IN4(\fadd_0_0_0_0_0/syncx_d2 [2]), .Q(n8360) );
  AO221X1 U882 ( .IN1(n8947), .IN2(n8364), .IN3(n14911), .IN4(n13956), .IN5(
        n8982), .Q(n12954) );
  AO22X1 U883 ( .IN1(n14910), .IN2(n13534), .IN3(n14421), .IN4(n13831), .Q(
        n8982) );
  AO22X1 U886 ( .IN1(\fadd_0_0_0_0_0/resultrounded [1]), .IN2(n14957), .IN3(
        n8958), .IN4(\fadd_0_0_0_0_0/syncx_d2 [1]), .Q(n8364) );
  AO221X1 U887 ( .IN1(n8947), .IN2(n8368), .IN3(n14911), .IN4(n13955), .IN5(
        n8984), .Q(n12955) );
  AO22X1 U888 ( .IN1(n14910), .IN2(n13523), .IN3(n14420), .IN4(n13830), .Q(
        n8984) );
  AO22X1 U891 ( .IN1(\fadd_0_0_0_0_0/resultrounded [0]), .IN2(n14957), .IN3(
        n8958), .IN4(\fadd_0_0_0_0_0/syncx_d2 [0]), .Q(n8368) );
  NAND4X0 U893 ( .IN1(n12146), .IN2(n12147), .IN3(n12148), .IN4(n13729), .QN(
        n8958) );
  AOI222X1 U899 ( .IN1(\U565/DATA1_11 ), .IN2(n14421), .IN3(n8989), .IN4(n8993), .IN5(n14911), .IN6(n13812), .QN(n8992) );
  NAND3X0 U902 ( .IN1(\fmul_0_0_0_0_0/expsigpostround [9]), .IN2(n14894), 
        .IN3(n11954), .QN(n8994) );
  OA222X1 U904 ( .IN1(n11952), .IN2(n8996), .IN3(n12696), .IN4(n8997), .IN5(
        n8998), .IN6(n8999), .Q(n8991) );
  AOI222X1 U906 ( .IN1(\U565/DATA1_10 ), .IN2(n14421), .IN3(n9002), .IN4(
        n11954), .IN5(n14911), .IN6(n13813), .QN(n9001) );
  OA21X1 U908 ( .IN1(n9003), .IN2(n13754), .IN3(n8989), .Q(n9002) );
  OA222X1 U911 ( .IN1(n11952), .IN2(n14765), .IN3(n11813), .IN4(n8997), .IN5(
        n14712), .IN6(n8999), .Q(n9000) );
  AOI222X1 U915 ( .IN1(\U565/DATA1_9 ), .IN2(n14421), .IN3(n14911), .IN4(
        n13811), .IN5(n8989), .IN6(\U565/DATA2_9 ), .QN(n9008) );
  OA222X1 U918 ( .IN1(n11952), .IN2(n9010), .IN3(n11812), .IN4(n8997), .IN5(
        n8523), .IN6(n8999), .Q(n9007) );
  OA222X1 U920 ( .IN1(n12332), .IN2(n9009), .IN3(n14713), .IN4(n8999), .IN5(
        n11952), .IN6(n14766), .Q(n9012) );
  AOI222X1 U923 ( .IN1(n14910), .IN2(n5986), .IN3(\U565/DATA2_8 ), .IN4(n8989), 
        .IN5(\U565/DATA1_8 ), .IN6(n14420), .QN(n9011) );
  OA222X1 U925 ( .IN1(n12334), .IN2(n9009), .IN3(n14714), .IN4(n8999), .IN5(
        n11952), .IN6(n14767), .Q(n9017) );
  AOI222X1 U928 ( .IN1(n14910), .IN2(n5985), .IN3(\U565/DATA2_7 ), .IN4(n8989), 
        .IN5(\U565/DATA1_7 ), .IN6(n14420), .QN(n9016) );
  OA222X1 U930 ( .IN1(n12336), .IN2(n9009), .IN3(n14715), .IN4(n8999), .IN5(
        n11952), .IN6(n14768), .Q(n9022) );
  AOI222X1 U933 ( .IN1(n14910), .IN2(n5984), .IN3(\U565/DATA2_6 ), .IN4(n8989), 
        .IN5(\U565/DATA1_6 ), .IN6(n14420), .QN(n9021) );
  OA222X1 U935 ( .IN1(n12338), .IN2(n9009), .IN3(n14716), .IN4(n8999), .IN5(
        n11952), .IN6(n14769), .Q(n9027) );
  AOI222X1 U938 ( .IN1(n14910), .IN2(n5983), .IN3(\U565/DATA2_5 ), .IN4(n8989), 
        .IN5(\U565/DATA1_5 ), .IN6(n14420), .QN(n9026) );
  OA222X1 U940 ( .IN1(n12340), .IN2(n9009), .IN3(n14717), .IN4(n8999), .IN5(
        n11952), .IN6(n14770), .Q(n9032) );
  AOI222X1 U943 ( .IN1(n14910), .IN2(n5982), .IN3(\U565/DATA2_4 ), .IN4(n8989), 
        .IN5(\U565/DATA1_4 ), .IN6(n14420), .QN(n9031) );
  OA222X1 U945 ( .IN1(n12342), .IN2(n9009), .IN3(n14718), .IN4(n8999), .IN5(
        n11952), .IN6(n14771), .Q(n9037) );
  AOI222X1 U948 ( .IN1(n14910), .IN2(n13713), .IN3(\U565/DATA2_3 ), .IN4(n8989), .IN5(\U565/DATA1_3 ), .IN6(n14420), .QN(n9036) );
  OA222X1 U950 ( .IN1(n12344), .IN2(n9009), .IN3(n14719), .IN4(n8999), .IN5(
        n11952), .IN6(n14772), .Q(n9042) );
  AOI222X1 U953 ( .IN1(n14910), .IN2(n13691), .IN3(\U565/DATA2_2 ), .IN4(n8989), .IN5(\U565/DATA1_2 ), .IN6(n14420), .QN(n9041) );
  OA222X1 U955 ( .IN1(n12346), .IN2(n9009), .IN3(n14720), .IN4(n8999), .IN5(
        n11952), .IN6(n14773), .Q(n9047) );
  AOI222X1 U958 ( .IN1(n14910), .IN2(n13670), .IN3(\U565/DATA2_1 ), .IN4(n8989), .IN5(\U565/DATA1_1 ), .IN6(n14420), .QN(n9046) );
  OA222X1 U960 ( .IN1(n12348), .IN2(n9009), .IN3(n14721), .IN4(n8999), .IN5(
        n11952), .IN6(n14774), .Q(n9052) );
  AOI222X1 U965 ( .IN1(n14910), .IN2(n13642), .IN3(\U565/DATA2_0 ), .IN4(n8989), .IN5(\U565/DATA1_0 ), .IN6(n14420), .QN(n9051) );
  AO221X1 U971 ( .IN1(n9058), .IN2(n14763), .IN3(n14417), .IN4(n13942), .IN5(
        n9060), .Q(n12968) );
  AO22X1 U972 ( .IN1(n9057), .IN2(n13514), .IN3(n9062), .IN4(n13817), .Q(n9060) );
  OA21X1 U976 ( .IN1(n14124), .IN2(n14764), .IN3(n12176), .Q(n8996) );
  AO221X1 U978 ( .IN1(n9058), .IN2(n8407), .IN3(n14417), .IN4(n13943), .IN5(
        n9066), .Q(n12969) );
  AO22X1 U979 ( .IN1(n9057), .IN2(n13505), .IN3(n9062), .IN4(n13818), .Q(n9066) );
  AO221X1 U982 ( .IN1(n9065), .IN2(n14124), .IN3(n9068), .IN4(n13725), .IN5(
        n9070), .Q(n8407) );
  NOR3X0 U985 ( .IN1(\fadd_0_0_0_0_4/resultrounded [10]), .IN2(n9068), .IN3(
        \fadd_0_0_0_0_4/zerofromclose_d1 ), .QN(n9065) );
  AO221X1 U986 ( .IN1(n14954), .IN2(n9058), .IN3(n14417), .IN4(n13941), .IN5(
        n9071), .Q(n12970) );
  AO22X1 U987 ( .IN1(n9057), .IN2(n13584), .IN3(n9062), .IN4(n13816), .Q(n9071) );
  AO22X1 U991 ( .IN1(n12179), .IN2(n14955), .IN3(n9074), .IN4(n9068), .Q(n9010) );
  NAND4X0 U993 ( .IN1(n12174), .IN2(n12175), .IN3(n9076), .IN4(n12176), .QN(
        n9075) );
  AO221X1 U996 ( .IN1(n9058), .IN2(n8380), .IN3(n14417), .IN4(n13952), .IN5(
        n9078), .Q(n12971) );
  AO22X1 U997 ( .IN1(n9057), .IN2(n5710), .IN3(n9062), .IN4(n13827), .Q(n9078)
         );
  AO22X1 U1000 ( .IN1(\fadd_0_0_0_0_4/resultrounded [8]), .IN2(n14955), .IN3(
        n9068), .IN4(\fadd_0_0_0_0_4/syncx_d2 [8]), .Q(n8380) );
  AO221X1 U1001 ( .IN1(n9058), .IN2(n8383), .IN3(n14417), .IN4(n13951), .IN5(
        n9080), .Q(n12972) );
  AO22X1 U1002 ( .IN1(n9057), .IN2(n5709), .IN3(n9062), .IN4(n13826), .Q(n9080) );
  AO22X1 U1005 ( .IN1(\fadd_0_0_0_0_4/resultrounded [7]), .IN2(n14955), .IN3(
        n9068), .IN4(\fadd_0_0_0_0_4/syncx_d2 [7]), .Q(n8383) );
  AO221X1 U1006 ( .IN1(n9058), .IN2(n8386), .IN3(n14417), .IN4(n13950), .IN5(
        n9082), .Q(n12973) );
  AO22X1 U1007 ( .IN1(n9057), .IN2(n5708), .IN3(n9062), .IN4(n13825), .Q(n9082) );
  AO22X1 U1010 ( .IN1(\fadd_0_0_0_0_4/resultrounded [6]), .IN2(n14955), .IN3(
        n9068), .IN4(\fadd_0_0_0_0_4/syncx_d2 [6]), .Q(n8386) );
  AO221X1 U1011 ( .IN1(n9058), .IN2(n8389), .IN3(n14417), .IN4(n13949), .IN5(
        n9084), .Q(n12974) );
  AO22X1 U1012 ( .IN1(n9057), .IN2(n5707), .IN3(n9062), .IN4(n13824), .Q(n9084) );
  AO22X1 U1015 ( .IN1(\fadd_0_0_0_0_4/resultrounded [5]), .IN2(n14955), .IN3(
        n9068), .IN4(\fadd_0_0_0_0_4/syncx_d2 [5]), .Q(n8389) );
  AO221X1 U1016 ( .IN1(n9058), .IN2(n8392), .IN3(n14417), .IN4(n13948), .IN5(
        n9086), .Q(n12975) );
  AO22X1 U1017 ( .IN1(n9057), .IN2(n5706), .IN3(n9062), .IN4(n13823), .Q(n9086) );
  AO22X1 U1020 ( .IN1(\fadd_0_0_0_0_4/resultrounded [4]), .IN2(n14955), .IN3(
        n9068), .IN4(\fadd_0_0_0_0_4/syncx_d2 [4]), .Q(n8392) );
  AO221X1 U1021 ( .IN1(n9058), .IN2(n8395), .IN3(n14417), .IN4(n13947), .IN5(
        n9088), .Q(n12976) );
  AO22X1 U1022 ( .IN1(n9057), .IN2(n13575), .IN3(n9062), .IN4(n13822), .Q(
        n9088) );
  AO22X1 U1025 ( .IN1(\fadd_0_0_0_0_4/resultrounded [3]), .IN2(n14955), .IN3(
        n9068), .IN4(\fadd_0_0_0_0_4/syncx_d2 [3]), .Q(n8395) );
  AO221X1 U1026 ( .IN1(n9058), .IN2(n8398), .IN3(n14417), .IN4(n13946), .IN5(
        n9090), .Q(n12977) );
  AO22X1 U1027 ( .IN1(n9057), .IN2(n13558), .IN3(n9062), .IN4(n13821), .Q(
        n9090) );
  AO22X1 U1030 ( .IN1(\fadd_0_0_0_0_4/resultrounded [2]), .IN2(n14955), .IN3(
        n9068), .IN4(\fadd_0_0_0_0_4/syncx_d2 [2]), .Q(n8398) );
  AO221X1 U1031 ( .IN1(n9058), .IN2(n8401), .IN3(n14417), .IN4(n13945), .IN5(
        n9092), .Q(n12978) );
  AO22X1 U1032 ( .IN1(n9057), .IN2(n13533), .IN3(n9062), .IN4(n13820), .Q(
        n9092) );
  AO22X1 U1035 ( .IN1(\fadd_0_0_0_0_4/resultrounded [1]), .IN2(n14955), .IN3(
        n9068), .IN4(\fadd_0_0_0_0_4/syncx_d2 [1]), .Q(n8401) );
  AO221X1 U1036 ( .IN1(n9058), .IN2(n8404), .IN3(n14417), .IN4(n13944), .IN5(
        n9094), .Q(n12979) );
  AO22X1 U1037 ( .IN1(n9057), .IN2(n13522), .IN3(n9062), .IN4(n13819), .Q(
        n9094) );
  AO22X1 U1040 ( .IN1(\fadd_0_0_0_0_4/resultrounded [0]), .IN2(n14955), .IN3(
        n9068), .IN4(\fadd_0_0_0_0_4/syncx_d2 [0]), .Q(n8404) );
  AO21X1 U1044 ( .IN1(n9096), .IN2(n8990), .IN3(n8988), .Q(n9058) );
  AO21X1 U1045 ( .IN1(n8764), .IN2(n9097), .IN3(n14184), .Q(n8988) );
  AO221X1 U1046 ( .IN1(n9057), .IN2(n13621), .IN3(n8449), .IN4(n14184), .IN5(
        n9099), .Q(n12980) );
  AO222X1 U1047 ( .IN1(n14417), .IN2(n13791), .IN3(n9096), .IN4(n9100), .IN5(
        \U341/DATA1_11 ), .IN6(n9062), .Q(n9099) );
  NAND3X0 U1049 ( .IN1(n14898), .IN2(n13747), .IN3(
        \fmul_0_0_0_0_4/expsigpostround [9]), .QN(n9102) );
  AO221X1 U1053 ( .IN1(n9057), .IN2(n13888), .IN3(n8446), .IN4(n14917), .IN5(
        n9106), .Q(n12981) );
  AO222X1 U1054 ( .IN1(n14418), .IN2(n13792), .IN3(n9107), .IN4(n9096), .IN5(
        \U341/DATA1_10 ), .IN6(n9062), .Q(n9106) );
  OA21X1 U1055 ( .IN1(n9108), .IN2(n11951), .IN3(n13747), .Q(n9107) );
  AO221X1 U1059 ( .IN1(n9057), .IN2(n13716), .IN3(n8416), .IN4(n14184), .IN5(
        n9110), .Q(n12982) );
  AO222X1 U1060 ( .IN1(\U341/DATA1_9 ), .IN2(n9062), .IN3(n14417), .IN4(n13779), .IN5(n9096), .IN6(\U341/DATA2_9 ), .Q(n9110) );
  AO221X1 U1062 ( .IN1(\U341/DATA2_8 ), .IN2(n9096), .IN3(n9057), .IN4(n5698), 
        .IN5(n9112), .Q(n12983) );
  AO222X1 U1063 ( .IN1(n14418), .IN2(n13810), .IN3(n8428), .IN4(n14917), .IN5(
        \U341/DATA1_8 ), .IN6(n9062), .Q(n9112) );
  AO221X1 U1065 ( .IN1(\U341/DATA2_7 ), .IN2(n9096), .IN3(n9057), .IN4(n5697), 
        .IN5(n9114), .Q(n12984) );
  AO222X1 U1066 ( .IN1(n14418), .IN2(n13809), .IN3(n8431), .IN4(n14917), .IN5(
        \U341/DATA1_7 ), .IN6(n9062), .Q(n9114) );
  AO221X1 U1068 ( .IN1(\U341/DATA2_6 ), .IN2(n9096), .IN3(n9057), .IN4(n5696), 
        .IN5(n9116), .Q(n12985) );
  AO222X1 U1069 ( .IN1(n14418), .IN2(n13808), .IN3(n8434), .IN4(n14917), .IN5(
        \U341/DATA1_6 ), .IN6(n9062), .Q(n9116) );
  AO221X1 U1071 ( .IN1(\U341/DATA2_5 ), .IN2(n9096), .IN3(n9057), .IN4(n5695), 
        .IN5(n9118), .Q(n12986) );
  AO222X1 U1072 ( .IN1(n14418), .IN2(n13807), .IN3(n8437), .IN4(n14917), .IN5(
        \U341/DATA1_5 ), .IN6(n9062), .Q(n9118) );
  AO221X1 U1074 ( .IN1(\U341/DATA2_4 ), .IN2(n9096), .IN3(n9057), .IN4(n5694), 
        .IN5(n9120), .Q(n12987) );
  AO222X1 U1075 ( .IN1(n14418), .IN2(n13806), .IN3(n8440), .IN4(n14184), .IN5(
        \U341/DATA1_4 ), .IN6(n9062), .Q(n9120) );
  AO221X1 U1077 ( .IN1(\U341/DATA2_3 ), .IN2(n9096), .IN3(n9057), .IN4(n13707), 
        .IN5(n9122), .Q(n12988) );
  AO222X1 U1078 ( .IN1(n14418), .IN2(n13805), .IN3(n8443), .IN4(n14917), .IN5(
        \U341/DATA1_3 ), .IN6(n9062), .Q(n9122) );
  AO221X1 U1080 ( .IN1(\U341/DATA2_2 ), .IN2(n9096), .IN3(n9057), .IN4(n13685), 
        .IN5(n9124), .Q(n12989) );
  AO222X1 U1081 ( .IN1(n14418), .IN2(n13804), .IN3(n8425), .IN4(n14917), .IN5(
        \U341/DATA1_2 ), .IN6(n9062), .Q(n9124) );
  AO221X1 U1083 ( .IN1(\U341/DATA2_1 ), .IN2(n9096), .IN3(n9057), .IN4(n13664), 
        .IN5(n9126), .Q(n12990) );
  AO222X1 U1084 ( .IN1(n14418), .IN2(n13803), .IN3(n8422), .IN4(n14917), .IN5(
        \U341/DATA1_1 ), .IN6(n9062), .Q(n9126) );
  AO221X1 U1086 ( .IN1(n13466), .IN2(n9096), .IN3(n9057), .IN4(n13636), .IN5(
        n9128), .Q(n12991) );
  AO222X1 U1087 ( .IN1(n14418), .IN2(n13802), .IN3(n8419), .IN4(n14184), .IN5(
        p___constant_11xf32_4[0]), .IN6(n9062), .Q(n9128) );
  AO221X1 U1095 ( .IN1(n14415), .IN2(n8449), .IN3(n14215), .IN4(n13929), .IN5(
        n9132), .Q(n12992) );
  AO22X1 U1096 ( .IN1(n14187), .IN2(n13859), .IN3(n14251), .IN4(n13508), .Q(
        n9132) );
  AO21X1 U1099 ( .IN1(\fadd_0_0_0_0_6/resultrounded [9]), .IN2(n9134), .IN3(
        n13777), .Q(n8449) );
  AO221X1 U1101 ( .IN1(n14415), .IN2(n8446), .IN3(n14215), .IN4(n13930), .IN5(
        n9136), .Q(n12993) );
  AO22X1 U1102 ( .IN1(n14263), .IN2(n13860), .IN3(n14251), .IN4(n13473), .Q(
        n9136) );
  AO221X1 U1105 ( .IN1(n9134), .IN2(n14816), .IN3(n9139), .IN4(n13728), .IN5(
        n9141), .Q(n8446) );
  NOR3X0 U1108 ( .IN1(\fadd_0_0_0_0_6/resultrounded [10]), .IN2(n9139), .IN3(
        \fadd_0_0_0_0_6/zerofromclose_d1 ), .QN(n9134) );
  AO221X1 U1109 ( .IN1(n14415), .IN2(n8416), .IN3(n14215), .IN4(n13940), .IN5(
        n9142), .Q(n12994) );
  OAI22X1 U1110 ( .IN1(n12828), .IN2(n12181), .IN3(n9130), .IN4(n11781), .QN(
        n9142) );
  AOI22X1 U1112 ( .IN1(n12182), .IN2(n14952), .IN3(n9144), .IN4(n9139), .QN(
        n8416) );
  NAND4X0 U1114 ( .IN1(n12209), .IN2(n13746), .IN3(n12207), .IN4(n9147), .QN(
        n9145) );
  AO221X1 U1117 ( .IN1(n14415), .IN2(n8428), .IN3(n14215), .IN4(n13936), .IN5(
        n9148), .Q(n12995) );
  AO22X1 U1118 ( .IN1(n14187), .IN2(n13866), .IN3(n14251), .IN4(n5566), .Q(
        n9148) );
  AO22X1 U1121 ( .IN1(\fadd_0_0_0_0_6/resultrounded [8]), .IN2(n14952), .IN3(
        n9139), .IN4(\fadd_0_0_0_0_6/syncx_d2 [8]), .Q(n8428) );
  AO221X1 U1122 ( .IN1(n14415), .IN2(n8431), .IN3(n14215), .IN4(n13935), .IN5(
        n9150), .Q(n12996) );
  AO22X1 U1123 ( .IN1(n14263), .IN2(n13865), .IN3(n14251), .IN4(n5565), .Q(
        n9150) );
  AO22X1 U1126 ( .IN1(\fadd_0_0_0_0_6/resultrounded [7]), .IN2(n14952), .IN3(
        n9139), .IN4(\fadd_0_0_0_0_6/syncx_d2 [7]), .Q(n8431) );
  AO221X1 U1127 ( .IN1(n14415), .IN2(n8434), .IN3(n14215), .IN4(n13934), .IN5(
        n9152), .Q(n12997) );
  AO22X1 U1128 ( .IN1(n14187), .IN2(n13864), .IN3(n14251), .IN4(n5564), .Q(
        n9152) );
  AO22X1 U1131 ( .IN1(\fadd_0_0_0_0_6/resultrounded [6]), .IN2(n14952), .IN3(
        n9139), .IN4(\fadd_0_0_0_0_6/syncx_d2 [6]), .Q(n8434) );
  AO221X1 U1132 ( .IN1(n14415), .IN2(n8437), .IN3(n14215), .IN4(n13933), .IN5(
        n9154), .Q(n12998) );
  AO22X1 U1133 ( .IN1(n14263), .IN2(n13863), .IN3(n14251), .IN4(n5563), .Q(
        n9154) );
  AO22X1 U1136 ( .IN1(\fadd_0_0_0_0_6/resultrounded [5]), .IN2(n14952), .IN3(
        n9139), .IN4(\fadd_0_0_0_0_6/syncx_d2 [5]), .Q(n8437) );
  AO221X1 U1137 ( .IN1(n14415), .IN2(n8440), .IN3(n14215), .IN4(n13932), .IN5(
        n9156), .Q(n12999) );
  AO22X1 U1138 ( .IN1(n14187), .IN2(n13862), .IN3(n14251), .IN4(n5562), .Q(
        n9156) );
  AO22X1 U1141 ( .IN1(\fadd_0_0_0_0_6/resultrounded [4]), .IN2(n14952), .IN3(
        n9139), .IN4(\fadd_0_0_0_0_6/syncx_d2 [4]), .Q(n8440) );
  AO221X1 U1142 ( .IN1(n14415), .IN2(n8443), .IN3(n14215), .IN4(n13931), .IN5(
        n9158), .Q(n13000) );
  AO22X1 U1143 ( .IN1(n14263), .IN2(n13861), .IN3(n14251), .IN4(n13496), .Q(
        n9158) );
  AO22X1 U1146 ( .IN1(\fadd_0_0_0_0_6/resultrounded [3]), .IN2(n14952), .IN3(
        n9139), .IN4(\fadd_0_0_0_0_6/syncx_d2 [3]), .Q(n8443) );
  AO221X1 U1147 ( .IN1(n14415), .IN2(n8425), .IN3(n14215), .IN4(n13937), .IN5(
        n9160), .Q(n13001) );
  AO22X1 U1148 ( .IN1(n14187), .IN2(n13867), .IN3(n14251), .IN4(n13494), .Q(
        n9160) );
  AO22X1 U1151 ( .IN1(\fadd_0_0_0_0_6/resultrounded [2]), .IN2(n14952), .IN3(
        n9139), .IN4(\fadd_0_0_0_0_6/syncx_d2 [2]), .Q(n8425) );
  AO221X1 U1152 ( .IN1(n14415), .IN2(n8422), .IN3(n14215), .IN4(n13938), .IN5(
        n9162), .Q(n13002) );
  AO22X1 U1153 ( .IN1(n14263), .IN2(n13868), .IN3(n14251), .IN4(n13481), .Q(
        n9162) );
  AO22X1 U1156 ( .IN1(\fadd_0_0_0_0_6/resultrounded [1]), .IN2(n14952), .IN3(
        n9139), .IN4(\fadd_0_0_0_0_6/syncx_d2 [1]), .Q(n8422) );
  AO221X1 U1157 ( .IN1(n14415), .IN2(n8419), .IN3(n14215), .IN4(n13939), .IN5(
        n9164), .Q(n13003) );
  AO22X1 U1158 ( .IN1(n14187), .IN2(n13869), .IN3(n14251), .IN4(n13479), .Q(
        n9164) );
  AO22X1 U1161 ( .IN1(\fadd_0_0_0_0_6/resultrounded [0]), .IN2(n14952), .IN3(
        n9139), .IN4(\fadd_0_0_0_0_6/syncx_d2 [0]), .Q(n8419) );
  NAND4X0 U1163 ( .IN1(n12207), .IN2(n12208), .IN3(n12209), .IN4(n13728), .QN(
        n9139) );
  AO221X1 U1165 ( .IN1(n9166), .IN2(n9167), .IN3(\U229/DATA1_11 ), .IN4(n14215), .IN5(n9168), .Q(n13004) );
  AO22X1 U1166 ( .IN1(n14263), .IN2(n13854), .IN3(n14251), .IN4(n13471), .Q(
        n9168) );
  NAND3X0 U1169 ( .IN1(n14900), .IN2(n13752), .IN3(
        \fmul_0_0_0_0_6/expsigpostround [9]), .QN(n9171) );
  AO221X1 U1172 ( .IN1(n9174), .IN2(n9166), .IN3(\U229/DATA1_10 ), .IN4(n14215), .IN5(n9175), .Q(n13005) );
  AO22X1 U1173 ( .IN1(n14187), .IN2(n13857), .IN3(n14251), .IN4(n13590), .Q(
        n9175) );
  OA21X1 U1175 ( .IN1(n9177), .IN2(n11949), .IN3(n13752), .Q(n9174) );
  AO221X1 U1178 ( .IN1(\U229/DATA1_9 ), .IN2(n14436), .IN3(n9166), .IN4(
        \U229/DATA2_9 ), .IN5(n9178), .Q(n13006) );
  OAI22X1 U1179 ( .IN1(n12828), .IN2(n12211), .IN3(n9130), .IN4(n11770), .QN(
        n9178) );
  AO221X1 U1180 ( .IN1(\U229/DATA1_8 ), .IN2(n14436), .IN3(\U229/DATA2_8 ), 
        .IN4(n9166), .IN5(n9179), .Q(n13007) );
  AO22X1 U1181 ( .IN1(n14263), .IN2(n13883), .IN3(n14251), .IN4(n5554), .Q(
        n9179) );
  AO221X1 U1183 ( .IN1(\U229/DATA1_7 ), .IN2(n14436), .IN3(\U229/DATA2_7 ), 
        .IN4(n9166), .IN5(n9181), .Q(n13008) );
  AO22X1 U1184 ( .IN1(n14187), .IN2(n13882), .IN3(n14251), .IN4(n5553), .Q(
        n9181) );
  AO221X1 U1186 ( .IN1(\U229/DATA1_6 ), .IN2(n14215), .IN3(\U229/DATA2_6 ), 
        .IN4(n9166), .IN5(n9183), .Q(n13009) );
  AO22X1 U1187 ( .IN1(n14263), .IN2(n13856), .IN3(n14251), .IN4(n5552), .Q(
        n9183) );
  AO221X1 U1189 ( .IN1(p___constant_11xf32_6[5]), .IN2(n14436), .IN3(n13459), 
        .IN4(n9166), .IN5(n9185), .Q(n13010) );
  AO22X1 U1190 ( .IN1(n14263), .IN2(n13881), .IN3(n14252), .IN4(n5551), .Q(
        n9185) );
  AO221X1 U1192 ( .IN1(p___constant_11xf32_6[4]), .IN2(n14215), .IN3(n13460), 
        .IN4(n9166), .IN5(n9187), .Q(n13011) );
  AO22X1 U1193 ( .IN1(n14187), .IN2(n13858), .IN3(n14252), .IN4(n5550), .Q(
        n9187) );
  AO221X1 U1195 ( .IN1(p___constant_11xf32_6[3]), .IN2(n14436), .IN3(n13461), 
        .IN4(n9166), .IN5(n9189), .Q(n13012) );
  AO22X1 U1196 ( .IN1(n14187), .IN2(n13880), .IN3(n14252), .IN4(n13578), .Q(
        n9189) );
  AO221X1 U1198 ( .IN1(p___constant_11xf32_6[2]), .IN2(n14215), .IN3(n13462), 
        .IN4(n9166), .IN5(n9191), .Q(n13013) );
  AO22X1 U1199 ( .IN1(n14263), .IN2(n13855), .IN3(n14252), .IN4(n13561), .Q(
        n9191) );
  AO221X1 U1201 ( .IN1(p___constant_11xf32_6[1]), .IN2(n14436), .IN3(n13463), 
        .IN4(n9166), .IN5(n9193), .Q(n13014) );
  AO22X1 U1202 ( .IN1(n14263), .IN2(n13879), .IN3(n14252), .IN4(n13536), .Q(
        n9193) );
  AO221X1 U1204 ( .IN1(p___constant_11xf32_6[0]), .IN2(n14215), .IN3(n13464), 
        .IN4(n9166), .IN5(n9195), .Q(n13015) );
  AO22X1 U1205 ( .IN1(n14187), .IN2(n13853), .IN3(n14252), .IN4(n13525), .Q(
        n9195) );
  AO222X1 U1207 ( .IN1(n14207), .IN2(n13512), .IN3(n14430), .IN4(n8482), .IN5(
        n14202), .IN6(n14005), .Q(n13016) );
  AO21X1 U1209 ( .IN1(\fadd_0_0_0_0_7/resultrounded [9]), .IN2(n9198), .IN3(
        n13773), .Q(n8482) );
  AO222X1 U1211 ( .IN1(n14213), .IN2(n13475), .IN3(n14430), .IN4(n8479), .IN5(
        n14203), .IN6(n14006), .Q(n13017) );
  AO221X1 U1213 ( .IN1(n9198), .IN2(n14837), .IN3(n9202), .IN4(n13734), .IN5(
        n9204), .Q(n8479) );
  NOR3X0 U1216 ( .IN1(\fadd_0_0_0_0_7/resultrounded [10]), .IN2(n9202), .IN3(
        \fadd_0_0_0_0_7/zerofromclose_d1 ), .QN(n9198) );
  AO222X1 U1217 ( .IN1(n14210), .IN2(n13582), .IN3(n14430), .IN4(n8452), .IN5(
        n14205), .IN6(n14015), .Q(n13018) );
  AOI22X1 U1219 ( .IN1(n12212), .IN2(n14950), .IN3(n9207), .IN4(n9202), .QN(
        n8452) );
  NAND4X0 U1221 ( .IN1(n12238), .IN2(n13744), .IN3(n12237), .IN4(n9210), .QN(
        n9208) );
  AO222X1 U1224 ( .IN1(n14213), .IN2(n5494), .IN3(n14430), .IN4(n8455), .IN5(
        n14260), .IN6(n14014), .Q(n13019) );
  AO22X1 U1226 ( .IN1(\fadd_0_0_0_0_7/resultrounded [8]), .IN2(n14950), .IN3(
        n9202), .IN4(\fadd_0_0_0_0_7/syncx_d2 [8]), .Q(n8455) );
  AO222X1 U1227 ( .IN1(n8766), .IN2(n5493), .IN3(n14430), .IN4(n8458), .IN5(
        n14261), .IN6(n14013), .Q(n13020) );
  AO22X1 U1229 ( .IN1(\fadd_0_0_0_0_7/resultrounded [7]), .IN2(n14950), .IN3(
        n9202), .IN4(\fadd_0_0_0_0_7/syncx_d2 [7]), .Q(n8458) );
  AO222X1 U1230 ( .IN1(n14211), .IN2(n5492), .IN3(n14430), .IN4(n8461), .IN5(
        n14201), .IN6(n14012), .Q(n13021) );
  AO22X1 U1232 ( .IN1(\fadd_0_0_0_0_7/resultrounded [6]), .IN2(n14950), .IN3(
        n9202), .IN4(\fadd_0_0_0_0_7/syncx_d2 [6]), .Q(n8461) );
  AO222X1 U1233 ( .IN1(n14210), .IN2(n5491), .IN3(n14430), .IN4(n8464), .IN5(
        n14259), .IN6(n14011), .Q(n13022) );
  AO22X1 U1235 ( .IN1(\fadd_0_0_0_0_7/resultrounded [5]), .IN2(n14950), .IN3(
        n9202), .IN4(\fadd_0_0_0_0_7/syncx_d2 [5]), .Q(n8464) );
  AO222X1 U1236 ( .IN1(n14208), .IN2(n5490), .IN3(n14430), .IN4(n8467), .IN5(
        n14204), .IN6(n14010), .Q(n13023) );
  AO22X1 U1238 ( .IN1(\fadd_0_0_0_0_7/resultrounded [4]), .IN2(n14950), .IN3(
        n9202), .IN4(\fadd_0_0_0_0_7/syncx_d2 [4]), .Q(n8467) );
  AO222X1 U1239 ( .IN1(n14207), .IN2(n13573), .IN3(n14430), .IN4(n8470), .IN5(
        n14205), .IN6(n14009), .Q(n13024) );
  AO22X1 U1241 ( .IN1(\fadd_0_0_0_0_7/resultrounded [3]), .IN2(n14950), .IN3(
        n9202), .IN4(\fadd_0_0_0_0_7/syncx_d2 [3]), .Q(n8470) );
  AO222X1 U1242 ( .IN1(n14212), .IN2(n13556), .IN3(n14430), .IN4(n8473), .IN5(
        n14204), .IN6(n14008), .Q(n13025) );
  AO22X1 U1244 ( .IN1(\fadd_0_0_0_0_7/resultrounded [2]), .IN2(n14950), .IN3(
        n9202), .IN4(\fadd_0_0_0_0_7/syncx_d2 [2]), .Q(n8473) );
  AO222X1 U1245 ( .IN1(n14212), .IN2(n13531), .IN3(n14430), .IN4(n8476), .IN5(
        n14202), .IN6(n14007), .Q(n13026) );
  AO22X1 U1247 ( .IN1(\fadd_0_0_0_0_7/resultrounded [1]), .IN2(n14950), .IN3(
        n9202), .IN4(\fadd_0_0_0_0_7/syncx_d2 [1]), .Q(n8476) );
  AO222X1 U1248 ( .IN1(n14214), .IN2(n13520), .IN3(n14430), .IN4(n8485), .IN5(
        n14206), .IN6(n14004), .Q(n13027) );
  AO22X1 U1250 ( .IN1(\fadd_0_0_0_0_7/resultrounded [0]), .IN2(n14950), .IN3(
        n9202), .IN4(\fadd_0_0_0_0_7/syncx_d2 [0]), .Q(n8485) );
  NAND4X0 U1252 ( .IN1(n12237), .IN2(n12238), .IN3(n12239), .IN4(n13734), .QN(
        n9202) );
  AO222X1 U1254 ( .IN1(n14213), .IN2(n13625), .IN3(n14422), .IN4(n9221), .IN5(
        \U173/DATA1_11 ), .IN6(n14206), .Q(n13028) );
  AO222X1 U1259 ( .IN1(n14214), .IN2(n13892), .IN3(n9227), .IN4(n14424), .IN5(
        \U173/DATA1_10 ), .IN6(n14916), .Q(n13029) );
  OA21X1 U1260 ( .IN1(n9228), .IN2(n11947), .IN3(n13769), .Q(n9227) );
  AO222X1 U1263 ( .IN1(n14214), .IN2(n13720), .IN3(n14422), .IN4(
        \U173/DATA2_9 ), .IN5(\U173/DATA1_9 ), .IN6(n14205), .Q(n13030) );
  AO222X1 U1264 ( .IN1(n14213), .IN2(n5482), .IN3(\U173/DATA2_8 ), .IN4(n14424), .IN5(\U173/DATA1_8 ), .IN6(n14204), .Q(n13031) );
  AO222X1 U1265 ( .IN1(n14209), .IN2(n5481), .IN3(\U173/DATA2_7 ), .IN4(n14424), .IN5(\U173/DATA1_7 ), .IN6(n14206), .Q(n13032) );
  AO222X1 U1266 ( .IN1(n14212), .IN2(n5480), .IN3(\U173/DATA2_6 ), .IN4(n14424), .IN5(\U173/DATA1_6 ), .IN6(n14261), .Q(n13033) );
  AO222X1 U1267 ( .IN1(n14207), .IN2(n5479), .IN3(\U173/DATA2_5 ), .IN4(n14424), .IN5(\U173/DATA1_5 ), .IN6(n14916), .Q(n13034) );
  AO222X1 U1268 ( .IN1(n14209), .IN2(n5478), .IN3(\U173/DATA2_4 ), .IN4(n14424), .IN5(\U173/DATA1_4 ), .IN6(n14203), .Q(n13035) );
  AO222X1 U1269 ( .IN1(n14207), .IN2(n13711), .IN3(\U173/DATA2_3 ), .IN4(
        n14425), .IN5(\U173/DATA1_3 ), .IN6(n14203), .Q(n13036) );
  AO222X1 U1270 ( .IN1(n14213), .IN2(n13689), .IN3(\U173/DATA2_2 ), .IN4(
        n14425), .IN5(\U173/DATA1_2 ), .IN6(n14183), .Q(n13037) );
  AO222X1 U1271 ( .IN1(n14211), .IN2(n13668), .IN3(n13457), .IN4(n14425), 
        .IN5(p___constant_11xf32_7[1]), .IN6(n14262), .Q(n13038) );
  AO222X1 U1272 ( .IN1(n14434), .IN2(n13640), .IN3(n13458), .IN4(n14425), 
        .IN5(p___constant_11xf32_7[0]), .IN6(n14261), .Q(n13039) );
  AO222X1 U1273 ( .IN1(n14433), .IN2(n13511), .IN3(n14431), .IN4(n8518), .IN5(
        n14260), .IN6(n13993), .Q(n13040) );
  AO21X1 U1275 ( .IN1(\fadd_0_0_0_0_5/resultrounded [9]), .IN2(n9240), .IN3(
        n13772), .Q(n8518) );
  AO222X1 U1277 ( .IN1(n14434), .IN2(n13503), .IN3(n14431), .IN4(n8515), .IN5(
        n14202), .IN6(n13994), .Q(n13041) );
  AO221X1 U1279 ( .IN1(n9240), .IN2(n14795), .IN3(n9244), .IN4(n13733), .IN5(
        n9246), .Q(n8515) );
  NOR3X0 U1282 ( .IN1(\fadd_0_0_0_0_5/resultrounded [10]), .IN2(n9244), .IN3(
        \fadd_0_0_0_0_5/zerofromclose_d1 ), .QN(n9240) );
  AO222X1 U1283 ( .IN1(n14212), .IN2(n13581), .IN3(n14431), .IN4(n8488), .IN5(
        n14260), .IN6(n14003), .Q(n13042) );
  AOI22X1 U1285 ( .IN1(n12242), .IN2(n14948), .IN3(n9249), .IN4(n9244), .QN(
        n8488) );
  NAND4X0 U1287 ( .IN1(n12268), .IN2(n13743), .IN3(n12267), .IN4(n9252), .QN(
        n9250) );
  AO222X1 U1290 ( .IN1(n8766), .IN2(n5638), .IN3(n14431), .IN4(n8491), .IN5(
        n14262), .IN6(n14002), .Q(n13043) );
  AO22X1 U1292 ( .IN1(\fadd_0_0_0_0_5/resultrounded [8]), .IN2(n14948), .IN3(
        n9244), .IN4(\fadd_0_0_0_0_5/syncx_d2 [8]), .Q(n8491) );
  AO222X1 U1293 ( .IN1(n14207), .IN2(n5637), .IN3(n14431), .IN4(n8494), .IN5(
        n14916), .IN6(n14001), .Q(n13044) );
  AO22X1 U1295 ( .IN1(\fadd_0_0_0_0_5/resultrounded [7]), .IN2(n14948), .IN3(
        n9244), .IN4(\fadd_0_0_0_0_5/syncx_d2 [7]), .Q(n8494) );
  AO222X1 U1296 ( .IN1(n14212), .IN2(n5636), .IN3(n14431), .IN4(n8497), .IN5(
        n14183), .IN6(n14000), .Q(n13045) );
  AO22X1 U1298 ( .IN1(\fadd_0_0_0_0_5/resultrounded [6]), .IN2(n14948), .IN3(
        n9244), .IN4(\fadd_0_0_0_0_5/syncx_d2 [6]), .Q(n8497) );
  AO222X1 U1299 ( .IN1(n14208), .IN2(n5635), .IN3(n14431), .IN4(n8500), .IN5(
        n14260), .IN6(n13999), .Q(n13046) );
  AO22X1 U1301 ( .IN1(\fadd_0_0_0_0_5/resultrounded [5]), .IN2(n14948), .IN3(
        n9244), .IN4(\fadd_0_0_0_0_5/syncx_d2 [5]), .Q(n8500) );
  AO222X1 U1302 ( .IN1(n14207), .IN2(n5634), .IN3(n14431), .IN4(n8503), .IN5(
        n14201), .IN6(n13998), .Q(n13047) );
  AO22X1 U1304 ( .IN1(\fadd_0_0_0_0_5/resultrounded [4]), .IN2(n14948), .IN3(
        n9244), .IN4(\fadd_0_0_0_0_5/syncx_d2 [4]), .Q(n8503) );
  AO222X1 U1305 ( .IN1(n14212), .IN2(n13572), .IN3(n14431), .IN4(n8506), .IN5(
        n14203), .IN6(n13997), .Q(n13048) );
  AO22X1 U1307 ( .IN1(\fadd_0_0_0_0_5/resultrounded [3]), .IN2(n14948), .IN3(
        n9244), .IN4(\fadd_0_0_0_0_5/syncx_d2 [3]), .Q(n8506) );
  AO222X1 U1308 ( .IN1(n14434), .IN2(n13555), .IN3(n14431), .IN4(n8509), .IN5(
        n14204), .IN6(n13996), .Q(n13049) );
  AO22X1 U1310 ( .IN1(\fadd_0_0_0_0_5/resultrounded [2]), .IN2(n14948), .IN3(
        n9244), .IN4(\fadd_0_0_0_0_5/syncx_d2 [2]), .Q(n8509) );
  AO222X1 U1311 ( .IN1(n14433), .IN2(n13530), .IN3(n14431), .IN4(n8512), .IN5(
        n14205), .IN6(n13995), .Q(n13050) );
  AO22X1 U1313 ( .IN1(\fadd_0_0_0_0_5/resultrounded [1]), .IN2(n14948), .IN3(
        n9244), .IN4(\fadd_0_0_0_0_5/syncx_d2 [1]), .Q(n8512) );
  AO222X1 U1314 ( .IN1(n14433), .IN2(n13519), .IN3(n14431), .IN4(n8521), .IN5(
        n14260), .IN6(n13992), .Q(n13051) );
  AO22X1 U1316 ( .IN1(\fadd_0_0_0_0_5/resultrounded [0]), .IN2(n14948), .IN3(
        n9244), .IN4(\fadd_0_0_0_0_5/syncx_d2 [0]), .Q(n8521) );
  NAND4X0 U1318 ( .IN1(n12267), .IN2(n12268), .IN3(n12269), .IN4(n13733), .QN(
        n9244) );
  AO222X1 U1320 ( .IN1(n14212), .IN2(n13624), .IN3(n14422), .IN4(n9263), .IN5(
        \U282/DATA1_11 ), .IN6(n14202), .Q(n13052) );
  AO222X1 U1325 ( .IN1(n8766), .IN2(n13891), .IN3(n9269), .IN4(n14425), .IN5(
        \U282/DATA1_10 ), .IN6(n14260), .Q(n13053) );
  OA21X1 U1326 ( .IN1(n9270), .IN2(n11945), .IN3(n13768), .Q(n9269) );
  AO222X1 U1329 ( .IN1(n14209), .IN2(n13719), .IN3(n14422), .IN4(
        \U282/DATA2_9 ), .IN5(\U282/DATA1_9 ), .IN6(n14206), .Q(n13054) );
  AO222X1 U1330 ( .IN1(n14210), .IN2(n5626), .IN3(\U282/DATA2_8 ), .IN4(n14425), .IN5(\U282/DATA1_8 ), .IN6(n14204), .Q(n13055) );
  AO222X1 U1331 ( .IN1(n14214), .IN2(n5625), .IN3(\U282/DATA2_7 ), .IN4(n14425), .IN5(\U282/DATA1_7 ), .IN6(n14205), .Q(n13056) );
  AO222X1 U1332 ( .IN1(n14213), .IN2(n5624), .IN3(\U282/DATA2_6 ), .IN4(n14425), .IN5(\U282/DATA1_6 ), .IN6(n14206), .Q(n13057) );
  AO222X1 U1333 ( .IN1(n14214), .IN2(n5623), .IN3(\U282/DATA2_5 ), .IN4(n14425), .IN5(\U282/DATA1_5 ), .IN6(n14261), .Q(n13058) );
  AO222X1 U1334 ( .IN1(n14209), .IN2(n5622), .IN3(\U282/DATA2_4 ), .IN4(n14425), .IN5(\U282/DATA1_4 ), .IN6(n14201), .Q(n13059) );
  AO222X1 U1335 ( .IN1(n14210), .IN2(n13710), .IN3(\U282/DATA2_3 ), .IN4(
        n14425), .IN5(\U282/DATA1_3 ), .IN6(n14202), .Q(n13060) );
  AO222X1 U1336 ( .IN1(n14211), .IN2(n13688), .IN3(\U282/DATA2_2 ), .IN4(
        n14425), .IN5(\U282/DATA1_2 ), .IN6(n14260), .Q(n13061) );
  AO222X1 U1337 ( .IN1(n14209), .IN2(n13667), .IN3(\U282/DATA2_1 ), .IN4(
        n14426), .IN5(\U282/DATA1_1 ), .IN6(n14204), .Q(n13062) );
  AO222X1 U1338 ( .IN1(n14211), .IN2(n13639), .IN3(n13465), .IN4(n14426), 
        .IN5(p___constant_11xf32_5[0]), .IN6(n14201), .Q(n13063) );
  AO221X1 U1339 ( .IN1(n14416), .IN2(n14710), .IN3(n14215), .IN4(n13918), 
        .IN5(n9281), .Q(n13064) );
  AO22X1 U1340 ( .IN1(n14187), .IN2(n13843), .IN3(n14252), .IN4(n13507), .Q(
        n9281) );
  OA21X1 U1344 ( .IN1(n14125), .IN2(n14711), .IN3(n12297), .Q(n8998) );
  AO221X1 U1346 ( .IN1(n14416), .IN2(n8551), .IN3(n14215), .IN4(n13919), .IN5(
        n9286), .Q(n13065) );
  AO22X1 U1347 ( .IN1(n14263), .IN2(n13844), .IN3(n14252), .IN4(n13472), .Q(
        n9286) );
  AO221X1 U1350 ( .IN1(n9285), .IN2(n14125), .IN3(n9288), .IN4(n13727), .IN5(
        n9290), .Q(n8551) );
  NOR3X0 U1353 ( .IN1(\fadd_0_0_0_0_2/resultrounded [10]), .IN2(n9288), .IN3(
        \fadd_0_0_0_0_2/zerofromclose_d1 ), .QN(n9285) );
  AO221X1 U1354 ( .IN1(n14416), .IN2(n14944), .IN3(n14215), .IN4(n13928), 
        .IN5(n9291), .Q(n13066) );
  OAI22X1 U1355 ( .IN1(n12828), .IN2(n12271), .IN3(n9130), .IN4(n11718), .QN(
        n9291) );
  AO22X1 U1358 ( .IN1(n12272), .IN2(n14945), .IN3(n9293), .IN4(n9288), .Q(
        n8523) );
  NAND4X0 U1360 ( .IN1(n12298), .IN2(n13738), .IN3(n12297), .IN4(n9296), .QN(
        n9294) );
  AO221X1 U1363 ( .IN1(n14416), .IN2(n8557), .IN3(n14215), .IN4(n13917), .IN5(
        n9297), .Q(n13067) );
  AO22X1 U1364 ( .IN1(n14187), .IN2(n13842), .IN3(n14252), .IN4(n5854), .Q(
        n9297) );
  AO22X1 U1367 ( .IN1(\fadd_0_0_0_0_2/resultrounded [8]), .IN2(n14945), .IN3(
        n9288), .IN4(\fadd_0_0_0_0_2/syncx_d2 [8]), .Q(n8557) );
  AO221X1 U1368 ( .IN1(n14416), .IN2(n8527), .IN3(n14215), .IN4(n13927), .IN5(
        n9299), .Q(n13068) );
  AO22X1 U1369 ( .IN1(n14263), .IN2(n13852), .IN3(n14252), .IN4(n5853), .Q(
        n9299) );
  AO22X1 U1372 ( .IN1(\fadd_0_0_0_0_2/resultrounded [7]), .IN2(n14945), .IN3(
        n9288), .IN4(\fadd_0_0_0_0_2/syncx_d2 [7]), .Q(n8527) );
  AO221X1 U1373 ( .IN1(n14416), .IN2(n8530), .IN3(n14215), .IN4(n13926), .IN5(
        n9301), .Q(n13069) );
  AO22X1 U1374 ( .IN1(n14187), .IN2(n13851), .IN3(n14252), .IN4(n5852), .Q(
        n9301) );
  AO22X1 U1377 ( .IN1(\fadd_0_0_0_0_2/resultrounded [6]), .IN2(n14945), .IN3(
        n9288), .IN4(\fadd_0_0_0_0_2/syncx_d2 [6]), .Q(n8530) );
  AO221X1 U1378 ( .IN1(n14416), .IN2(n8533), .IN3(n14215), .IN4(n13925), .IN5(
        n9303), .Q(n13070) );
  AO22X1 U1379 ( .IN1(n14263), .IN2(n13850), .IN3(n14252), .IN4(n5851), .Q(
        n9303) );
  AO22X1 U1382 ( .IN1(\fadd_0_0_0_0_2/resultrounded [5]), .IN2(n14945), .IN3(
        n9288), .IN4(\fadd_0_0_0_0_2/syncx_d2 [5]), .Q(n8533) );
  AO221X1 U1383 ( .IN1(n14416), .IN2(n8536), .IN3(n14215), .IN4(n13924), .IN5(
        n9305), .Q(n13071) );
  AO22X1 U1384 ( .IN1(n14187), .IN2(n13849), .IN3(n14252), .IN4(n5850), .Q(
        n9305) );
  AO22X1 U1387 ( .IN1(\fadd_0_0_0_0_2/resultrounded [4]), .IN2(n14945), .IN3(
        n9288), .IN4(\fadd_0_0_0_0_2/syncx_d2 [4]), .Q(n8536) );
  AO221X1 U1388 ( .IN1(n14416), .IN2(n8539), .IN3(n14215), .IN4(n13923), .IN5(
        n9307), .Q(n13072) );
  AO22X1 U1389 ( .IN1(n14263), .IN2(n13848), .IN3(n14252), .IN4(n13495), .Q(
        n9307) );
  AO22X1 U1392 ( .IN1(\fadd_0_0_0_0_2/resultrounded [3]), .IN2(n14945), .IN3(
        n9288), .IN4(\fadd_0_0_0_0_2/syncx_d2 [3]), .Q(n8539) );
  AO221X1 U1393 ( .IN1(n14416), .IN2(n8542), .IN3(n14215), .IN4(n13922), .IN5(
        n9309), .Q(n13073) );
  AO22X1 U1394 ( .IN1(n14263), .IN2(n13847), .IN3(n14252), .IN4(n13493), .Q(
        n9309) );
  AO22X1 U1397 ( .IN1(\fadd_0_0_0_0_2/resultrounded [2]), .IN2(n14945), .IN3(
        n9288), .IN4(\fadd_0_0_0_0_2/syncx_d2 [2]), .Q(n8542) );
  AO221X1 U1398 ( .IN1(n14416), .IN2(n8545), .IN3(n14215), .IN4(n13921), .IN5(
        n9311), .Q(n13074) );
  AO22X1 U1399 ( .IN1(n14263), .IN2(n13846), .IN3(n14252), .IN4(n13480), .Q(
        n9311) );
  AO22X1 U1402 ( .IN1(\fadd_0_0_0_0_2/resultrounded [1]), .IN2(n14945), .IN3(
        n9288), .IN4(\fadd_0_0_0_0_2/syncx_d2 [1]), .Q(n8545) );
  AO221X1 U1403 ( .IN1(n14416), .IN2(n8548), .IN3(n14215), .IN4(n13920), .IN5(
        n9313), .Q(n13075) );
  AO22X1 U1404 ( .IN1(n14187), .IN2(n13845), .IN3(n14252), .IN4(n13478), .Q(
        n9313) );
  AO22X1 U1407 ( .IN1(\fadd_0_0_0_0_2/resultrounded [0]), .IN2(n14945), .IN3(
        n9288), .IN4(\fadd_0_0_0_0_2/syncx_d2 [0]), .Q(n8548) );
  AO221X1 U1412 ( .IN1(n9166), .IN2(n9315), .IN3(\U450/DATA1_11 ), .IN4(n14215), .IN5(n9316), .Q(n13076) );
  AO22X1 U1413 ( .IN1(n14187), .IN2(n13840), .IN3(n14253), .IN4(n13470), .Q(
        n9316) );
  NAND3X0 U1416 ( .IN1(n14896), .IN2(n13751), .IN3(
        \fmul_0_0_0_0_2/expsigpostround [9]), .QN(n9319) );
  AO221X1 U1419 ( .IN1(n9322), .IN2(n9166), .IN3(\U450/DATA1_10 ), .IN4(n14215), .IN5(n9323), .Q(n13077) );
  AO22X1 U1420 ( .IN1(n14187), .IN2(n13841), .IN3(n14253), .IN4(n13589), .Q(
        n9323) );
  OA21X1 U1422 ( .IN1(n9325), .IN2(n11943), .IN3(n13751), .Q(n9322) );
  AO221X1 U1425 ( .IN1(\U450/DATA1_9 ), .IN2(n14436), .IN3(n9166), .IN4(
        \U450/DATA2_9 ), .IN5(n9326), .Q(n13078) );
  OAI22X1 U1426 ( .IN1(n12828), .IN2(n12324), .IN3(n9130), .IN4(n11707), .QN(
        n9326) );
  AO221X1 U1427 ( .IN1(\U450/DATA1_8 ), .IN2(n14436), .IN3(\U450/DATA2_8 ), 
        .IN4(n9166), .IN5(n9327), .Q(n13079) );
  AO22X1 U1428 ( .IN1(n14263), .IN2(n13878), .IN3(n14253), .IN4(n5842), .Q(
        n9327) );
  AO221X1 U1430 ( .IN1(\U450/DATA1_7 ), .IN2(n14436), .IN3(\U450/DATA2_7 ), 
        .IN4(n9166), .IN5(n9329), .Q(n13080) );
  AO22X1 U1431 ( .IN1(n14263), .IN2(n13877), .IN3(n14253), .IN4(n5841), .Q(
        n9329) );
  AO221X1 U1433 ( .IN1(\U450/DATA1_6 ), .IN2(n14436), .IN3(\U450/DATA2_6 ), 
        .IN4(n9166), .IN5(n9331), .Q(n13081) );
  AO22X1 U1434 ( .IN1(n14263), .IN2(n13876), .IN3(n14253), .IN4(n5840), .Q(
        n9331) );
  AO221X1 U1436 ( .IN1(\U450/DATA1_5 ), .IN2(n14436), .IN3(\U450/DATA2_5 ), 
        .IN4(n9166), .IN5(n9333), .Q(n13082) );
  AO22X1 U1437 ( .IN1(n14187), .IN2(n13875), .IN3(n14253), .IN4(n5839), .Q(
        n9333) );
  AO221X1 U1439 ( .IN1(\U450/DATA1_4 ), .IN2(n14436), .IN3(\U450/DATA2_4 ), 
        .IN4(n9166), .IN5(n9335), .Q(n13083) );
  AO22X1 U1440 ( .IN1(n14187), .IN2(n13874), .IN3(n14253), .IN4(n5838), .Q(
        n9335) );
  AO221X1 U1442 ( .IN1(\U450/DATA1_3 ), .IN2(n14436), .IN3(\U450/DATA2_3 ), 
        .IN4(n9166), .IN5(n9337), .Q(n13084) );
  AO22X1 U1443 ( .IN1(n14187), .IN2(n13873), .IN3(n14253), .IN4(n13577), .Q(
        n9337) );
  AO221X1 U1445 ( .IN1(\U450/DATA1_2 ), .IN2(n14436), .IN3(\U450/DATA2_2 ), 
        .IN4(n9166), .IN5(n9339), .Q(n13085) );
  AO22X1 U1446 ( .IN1(n14187), .IN2(n13872), .IN3(n14253), .IN4(n13560), .Q(
        n9339) );
  AO221X1 U1448 ( .IN1(\U450/DATA1_1 ), .IN2(n14436), .IN3(\U450/DATA2_1 ), 
        .IN4(n9166), .IN5(n9341), .Q(n13086) );
  AO22X1 U1449 ( .IN1(n14263), .IN2(n13871), .IN3(n14253), .IN4(n13535), .Q(
        n9341) );
  AO221X1 U1451 ( .IN1(\U450/DATA1_0 ), .IN2(n14436), .IN3(\U450/DATA2_0 ), 
        .IN4(n9166), .IN5(n9343), .Q(n13087) );
  AO22X1 U1452 ( .IN1(n14263), .IN2(n13870), .IN3(n14253), .IN4(n13524), .Q(
        n9343) );
  AO222X1 U1460 ( .IN1(n14433), .IN2(n13510), .IN3(n14432), .IN4(n8590), .IN5(
        n14261), .IN6(n13981), .Q(n13088) );
  AO21X1 U1462 ( .IN1(\fadd_0_0_0_0_3/resultrounded [9]), .IN2(n9346), .IN3(
        n13775), .Q(n8590) );
  AO222X1 U1464 ( .IN1(n14213), .IN2(n13474), .IN3(n14432), .IN4(n8587), .IN5(
        n14204), .IN6(n13982), .Q(n13089) );
  AO221X1 U1466 ( .IN1(n9346), .IN2(n14742), .IN3(n9350), .IN4(n13731), .IN5(
        n9352), .Q(n8587) );
  NOR3X0 U1469 ( .IN1(\fadd_0_0_0_0_3/resultrounded [10]), .IN2(n9350), .IN3(
        \fadd_0_0_0_0_3/zerofromclose_d1 ), .QN(n9346) );
  AO222X1 U1470 ( .IN1(n14209), .IN2(n13580), .IN3(n14432), .IN4(n8593), .IN5(
        n14201), .IN6(n13980), .Q(n13090) );
  AOI22X1 U1472 ( .IN1(n12330), .IN2(n14943), .IN3(n9355), .IN4(n9350), .QN(
        n8593) );
  NAND4X0 U1474 ( .IN1(n12325), .IN2(n12326), .IN3(n9357), .IN4(n12327), .QN(
        n9356) );
  AO222X1 U1477 ( .IN1(n8766), .IN2(n5782), .IN3(n14432), .IN4(n8560), .IN5(
        n14201), .IN6(n13991), .Q(n13091) );
  AO22X1 U1479 ( .IN1(\fadd_0_0_0_0_3/resultrounded [8]), .IN2(n14943), .IN3(
        n9350), .IN4(\fadd_0_0_0_0_3/syncx_d2 [8]), .Q(n8560) );
  AO222X1 U1480 ( .IN1(n14214), .IN2(n5781), .IN3(n14432), .IN4(n8563), .IN5(
        n14206), .IN6(n13990), .Q(n13092) );
  AO22X1 U1482 ( .IN1(\fadd_0_0_0_0_3/resultrounded [7]), .IN2(n14943), .IN3(
        n9350), .IN4(\fadd_0_0_0_0_3/syncx_d2 [7]), .Q(n8563) );
  AO222X1 U1483 ( .IN1(n14213), .IN2(n5780), .IN3(n14432), .IN4(n8566), .IN5(
        n14259), .IN6(n13989), .Q(n13093) );
  AO22X1 U1485 ( .IN1(\fadd_0_0_0_0_3/resultrounded [6]), .IN2(n14943), .IN3(
        n9350), .IN4(\fadd_0_0_0_0_3/syncx_d2 [6]), .Q(n8566) );
  AO222X1 U1486 ( .IN1(n14210), .IN2(n5779), .IN3(n14432), .IN4(n8569), .IN5(
        n14259), .IN6(n13988), .Q(n13094) );
  AO22X1 U1488 ( .IN1(\fadd_0_0_0_0_3/resultrounded [5]), .IN2(n14943), .IN3(
        n9350), .IN4(\fadd_0_0_0_0_3/syncx_d2 [5]), .Q(n8569) );
  AO222X1 U1489 ( .IN1(n14211), .IN2(n5778), .IN3(n14432), .IN4(n8572), .IN5(
        n14206), .IN6(n13987), .Q(n13095) );
  AO22X1 U1491 ( .IN1(\fadd_0_0_0_0_3/resultrounded [4]), .IN2(n14943), .IN3(
        n9350), .IN4(\fadd_0_0_0_0_3/syncx_d2 [4]), .Q(n8572) );
  AO222X1 U1492 ( .IN1(n14208), .IN2(n13571), .IN3(n14432), .IN4(n8575), .IN5(
        n14261), .IN6(n13986), .Q(n13096) );
  AO22X1 U1494 ( .IN1(\fadd_0_0_0_0_3/resultrounded [3]), .IN2(n14943), .IN3(
        n9350), .IN4(\fadd_0_0_0_0_3/syncx_d2 [3]), .Q(n8575) );
  AO222X1 U1495 ( .IN1(n14208), .IN2(n13554), .IN3(n14432), .IN4(n8578), .IN5(
        n14203), .IN6(n13985), .Q(n13097) );
  AO22X1 U1497 ( .IN1(\fadd_0_0_0_0_3/resultrounded [2]), .IN2(n14943), .IN3(
        n9350), .IN4(\fadd_0_0_0_0_3/syncx_d2 [2]), .Q(n8578) );
  AO222X1 U1498 ( .IN1(n14434), .IN2(n13529), .IN3(n14432), .IN4(n8581), .IN5(
        n14203), .IN6(n13984), .Q(n13098) );
  AO22X1 U1500 ( .IN1(\fadd_0_0_0_0_3/resultrounded [1]), .IN2(n14943), .IN3(
        n9350), .IN4(\fadd_0_0_0_0_3/syncx_d2 [1]), .Q(n8581) );
  AO222X1 U1501 ( .IN1(n14433), .IN2(n13518), .IN3(n14432), .IN4(n8584), .IN5(
        n14205), .IN6(n13983), .Q(n13099) );
  AO22X1 U1503 ( .IN1(\fadd_0_0_0_0_3/resultrounded [0]), .IN2(n14943), .IN3(
        n9350), .IN4(\fadd_0_0_0_0_3/syncx_d2 [0]), .Q(n8584) );
  AO222X1 U1507 ( .IN1(n14208), .IN2(n13623), .IN3(n14422), .IN4(n9369), .IN5(
        \U394/DATA1_11 ), .IN6(n14262), .Q(n13100) );
  AO222X1 U1512 ( .IN1(n14433), .IN2(n13890), .IN3(n9375), .IN4(n14426), .IN5(
        \U394/DATA1_10 ), .IN6(n14202), .Q(n13101) );
  OA21X1 U1513 ( .IN1(n9376), .IN2(n11941), .IN3(n13767), .Q(n9375) );
  AO222X1 U1516 ( .IN1(n14211), .IN2(n13718), .IN3(n14422), .IN4(
        \U394/DATA2_9 ), .IN5(\U394/DATA1_9 ), .IN6(n14203), .Q(n13102) );
  AO222X1 U1517 ( .IN1(n8766), .IN2(n5770), .IN3(\U394/DATA2_8 ), .IN4(n14426), 
        .IN5(\U394/DATA1_8 ), .IN6(n14183), .Q(n13103) );
  AO222X1 U1518 ( .IN1(n14434), .IN2(n5769), .IN3(\U394/DATA2_7 ), .IN4(n14426), .IN5(\U394/DATA1_7 ), .IN6(n14205), .Q(n13104) );
  AO222X1 U1519 ( .IN1(n14433), .IN2(n5768), .IN3(\U394/DATA2_6 ), .IN4(n14426), .IN5(\U394/DATA1_6 ), .IN6(n14206), .Q(n13105) );
  AO222X1 U1520 ( .IN1(n14209), .IN2(n5767), .IN3(\U394/DATA2_5 ), .IN4(n14426), .IN5(\U394/DATA1_5 ), .IN6(n14202), .Q(n13106) );
  AO222X1 U1521 ( .IN1(n14207), .IN2(n5766), .IN3(\U394/DATA2_4 ), .IN4(n14426), .IN5(\U394/DATA1_4 ), .IN6(n14205), .Q(n13107) );
  AO222X1 U1522 ( .IN1(n14214), .IN2(n13709), .IN3(\U394/DATA2_3 ), .IN4(
        n14426), .IN5(\U394/DATA1_3 ), .IN6(n14205), .Q(n13108) );
  AO222X1 U1523 ( .IN1(n14433), .IN2(n13687), .IN3(\U394/DATA2_2 ), .IN4(
        n14426), .IN5(\U394/DATA1_2 ), .IN6(n14201), .Q(n13109) );
  AO222X1 U1524 ( .IN1(n14211), .IN2(n13666), .IN3(\U394/DATA2_1 ), .IN4(
        n14426), .IN5(\U394/DATA1_1 ), .IN6(n14259), .Q(n13110) );
  AO222X1 U1525 ( .IN1(n14210), .IN2(n13638), .IN3(\U394/DATA2_0 ), .IN4(
        n14426), .IN5(\U394/DATA1_0 ), .IN6(n14262), .Q(n13111) );
  AO222X1 U1526 ( .IN1(n14213), .IN2(n13509), .IN3(n14431), .IN4(n8626), .IN5(
        n14203), .IN6(n13969), .Q(n13112) );
  AO21X1 U1528 ( .IN1(\fadd_0_0_0_0_1/resultrounded [9]), .IN2(n9388), .IN3(
        n13774), .Q(n8626) );
  AO222X1 U1530 ( .IN1(n14210), .IN2(n13502), .IN3(n8768), .IN4(n8623), .IN5(
        n14201), .IN6(n13970), .Q(n13113) );
  AO221X1 U1532 ( .IN1(n9388), .IN2(n14689), .IN3(n9392), .IN4(n13730), .IN5(
        n9394), .Q(n8623) );
  NOR3X0 U1535 ( .IN1(\fadd_0_0_0_0_1/resultrounded [10]), .IN2(n9392), .IN3(
        \fadd_0_0_0_0_1/zerofromclose_d1 ), .QN(n9388) );
  AO222X1 U1536 ( .IN1(n14209), .IN2(n13579), .IN3(n14430), .IN4(n8629), .IN5(
        n14202), .IN6(n13968), .Q(n13114) );
  AOI22X1 U1538 ( .IN1(n12362), .IN2(n14941), .IN3(n9397), .IN4(n9392), .QN(
        n8629) );
  NAND4X0 U1540 ( .IN1(n12357), .IN2(n12358), .IN3(n9399), .IN4(n12359), .QN(
        n9398) );
  AO222X1 U1543 ( .IN1(n14207), .IN2(n5926), .IN3(n8768), .IN4(n8596), .IN5(
        n14205), .IN6(n13979), .Q(n13115) );
  AO22X1 U1545 ( .IN1(\fadd_0_0_0_0_1/resultrounded [8]), .IN2(n14941), .IN3(
        n9392), .IN4(\fadd_0_0_0_0_1/syncx_d2 [8]), .Q(n8596) );
  AO222X1 U1546 ( .IN1(n14211), .IN2(n5925), .IN3(n14429), .IN4(n8599), .IN5(
        n14202), .IN6(n13978), .Q(n13116) );
  AO22X1 U1548 ( .IN1(\fadd_0_0_0_0_1/resultrounded [7]), .IN2(n14941), .IN3(
        n9392), .IN4(\fadd_0_0_0_0_1/syncx_d2 [7]), .Q(n8599) );
  AO222X1 U1549 ( .IN1(n14210), .IN2(n5924), .IN3(n14432), .IN4(n8602), .IN5(
        n14202), .IN6(n13977), .Q(n13117) );
  AO22X1 U1551 ( .IN1(\fadd_0_0_0_0_1/resultrounded [6]), .IN2(n14941), .IN3(
        n9392), .IN4(\fadd_0_0_0_0_1/syncx_d2 [6]), .Q(n8602) );
  AO222X1 U1552 ( .IN1(n14208), .IN2(n5923), .IN3(n8768), .IN4(n8605), .IN5(
        n14206), .IN6(n13976), .Q(n13118) );
  AO22X1 U1554 ( .IN1(\fadd_0_0_0_0_1/resultrounded [5]), .IN2(n14941), .IN3(
        n9392), .IN4(\fadd_0_0_0_0_1/syncx_d2 [5]), .Q(n8605) );
  AO222X1 U1555 ( .IN1(n14207), .IN2(n5922), .IN3(n8768), .IN4(n8608), .IN5(
        n14206), .IN6(n13975), .Q(n13119) );
  AO22X1 U1557 ( .IN1(\fadd_0_0_0_0_1/resultrounded [4]), .IN2(n14941), .IN3(
        n9392), .IN4(\fadd_0_0_0_0_1/syncx_d2 [4]), .Q(n8608) );
  AO222X1 U1558 ( .IN1(n14212), .IN2(n13570), .IN3(n8768), .IN4(n8611), .IN5(
        n14204), .IN6(n13974), .Q(n13120) );
  AO22X1 U1560 ( .IN1(\fadd_0_0_0_0_1/resultrounded [3]), .IN2(n14941), .IN3(
        n9392), .IN4(\fadd_0_0_0_0_1/syncx_d2 [3]), .Q(n8611) );
  AO222X1 U1561 ( .IN1(n14207), .IN2(n13553), .IN3(n8768), .IN4(n8614), .IN5(
        n14259), .IN6(n13973), .Q(n13121) );
  AO22X1 U1563 ( .IN1(\fadd_0_0_0_0_1/resultrounded [2]), .IN2(n14941), .IN3(
        n9392), .IN4(\fadd_0_0_0_0_1/syncx_d2 [2]), .Q(n8614) );
  AO222X1 U1564 ( .IN1(n14434), .IN2(n13528), .IN3(n14428), .IN4(n8617), .IN5(
        n14205), .IN6(n13972), .Q(n13122) );
  AO22X1 U1566 ( .IN1(\fadd_0_0_0_0_1/resultrounded [1]), .IN2(n14941), .IN3(
        n9392), .IN4(\fadd_0_0_0_0_1/syncx_d2 [1]), .Q(n8617) );
  AO222X1 U1567 ( .IN1(n14210), .IN2(n13517), .IN3(n8768), .IN4(n8620), .IN5(
        n14204), .IN6(n13971), .Q(n13123) );
  AO22X1 U1569 ( .IN1(\fadd_0_0_0_0_1/resultrounded [0]), .IN2(n14941), .IN3(
        n9392), .IN4(\fadd_0_0_0_0_1/syncx_d2 [0]), .Q(n8620) );
  AND2X1 U1573 ( .IN1(n14427), .IN2(n14912), .Q(n8768) );
  AO222X1 U1575 ( .IN1(n8766), .IN2(n13622), .IN3(n14422), .IN4(n9412), .IN5(
        \U503/DATA1_11 ), .IN6(n14203), .Q(n13124) );
  AO222X1 U1580 ( .IN1(n14434), .IN2(n13889), .IN3(n9418), .IN4(n14426), .IN5(
        \U503/DATA1_10 ), .IN6(n14203), .Q(n13125) );
  OA21X1 U1581 ( .IN1(n9419), .IN2(n11939), .IN3(n13766), .Q(n9418) );
  AO222X1 U1584 ( .IN1(n14433), .IN2(n13717), .IN3(n14422), .IN4(
        \U503/DATA2_9 ), .IN5(\U503/DATA1_9 ), .IN6(n14201), .Q(n13126) );
  AO222X1 U1585 ( .IN1(n14210), .IN2(n5914), .IN3(\U503/DATA2_8 ), .IN4(n14427), .IN5(\U503/DATA1_8 ), .IN6(n14205), .Q(n13127) );
  AO222X1 U1586 ( .IN1(n14208), .IN2(n5913), .IN3(\U503/DATA2_7 ), .IN4(n14427), .IN5(\U503/DATA1_7 ), .IN6(n14204), .Q(n13128) );
  AO222X1 U1587 ( .IN1(n8766), .IN2(n5912), .IN3(\U503/DATA2_6 ), .IN4(n14427), 
        .IN5(\U503/DATA1_6 ), .IN6(n14202), .Q(n13129) );
  AO222X1 U1588 ( .IN1(n14214), .IN2(n5911), .IN3(\U503/DATA2_5 ), .IN4(n14427), .IN5(\U503/DATA1_5 ), .IN6(n14204), .Q(n13130) );
  AO222X1 U1589 ( .IN1(n14208), .IN2(n5910), .IN3(\U503/DATA2_4 ), .IN4(n14427), .IN5(\U503/DATA1_4 ), .IN6(n14261), .Q(n13131) );
  AO222X1 U1590 ( .IN1(n14434), .IN2(n13708), .IN3(\U503/DATA2_3 ), .IN4(
        n14427), .IN5(\U503/DATA1_3 ), .IN6(n14262), .Q(n13132) );
  AO222X1 U1591 ( .IN1(n14212), .IN2(n13686), .IN3(\U503/DATA2_2 ), .IN4(
        n14427), .IN5(\U503/DATA1_2 ), .IN6(n14916), .Q(n13133) );
  AO222X1 U1592 ( .IN1(n14214), .IN2(n13665), .IN3(\U503/DATA2_1 ), .IN4(
        n14427), .IN5(\U503/DATA1_1 ), .IN6(n14183), .Q(n13134) );
  AO222X1 U1593 ( .IN1(n14213), .IN2(n13637), .IN3(\U503/DATA2_0 ), .IN4(
        n14423), .IN5(\U503/DATA1_0 ), .IN6(n14259), .Q(n13135) );
  AND3X1 U1596 ( .IN1(n9410), .IN2(n12829), .IN3(n11937), .Q(n8766) );
  OR2X1 U1598 ( .IN1(n11935), .IN2(n11936), .Q(n9097) );
  NAND4X0 U1599 ( .IN1(n11929), .IN2(n11930), .IN3(n9430), .IN4(n9431), .QN(
        n8990) );
  AND4X1 U1600 ( .IN1(n13476), .IN2(n13631), .IN3(n11934), .IN4(n11933), .Q(
        n9431) );
  AND2X1 U1601 ( .IN1(n11932), .IN2(n11931), .Q(n9430) );
  AO221X1 U1603 ( .IN1(n14235), .IN2(n13916), .IN3(\U10/DATA1_11 ), .IN4(
        n14197), .IN5(n9439), .Q(n13137) );
  AO222X1 U1604 ( .IN1(\U15/DATA1_11 ), .IN2(n14410), .IN3(n14397), .IN4(n9442), .IN5(\U20/DATA1_11 ), .IN6(n14386), .Q(n9439) );
  OR2X1 U1605 ( .IN1(n9444), .IN2(n9445), .Q(n9442) );
  AO221X1 U1606 ( .IN1(\U50/DATA1_11 ), .IN2(n14385), .IN3(\U55/DATA1_11 ), 
        .IN4(n14373), .IN5(n9448), .Q(n9445) );
  AO22X1 U1607 ( .IN1(\U25/DATA1_11 ), .IN2(n14189), .IN3(\U55/DATA2_11 ), 
        .IN4(n14360), .Q(n9448) );
  AO221X1 U1608 ( .IN1(\U30/DATA1_11 ), .IN2(n14354), .IN3(\U45/DATA1_11 ), 
        .IN4(n14343), .IN5(n9453), .Q(n9444) );
  AO22X1 U1609 ( .IN1(\U35/DATA1_11 ), .IN2(n14333), .IN3(\U40/DATA1_11 ), 
        .IN4(n14322), .Q(n9453) );
  AO221X1 U1611 ( .IN1(n14235), .IN2(n13607), .IN3(\U10/DATA1_10 ), .IN4(
        n14196), .IN5(n9457), .Q(n13138) );
  AO222X1 U1612 ( .IN1(p___constant_11x11xf32_10_9[10]), .IN2(n14407), .IN3(
        n14397), .IN4(n9458), .IN5(\U20/DATA1_10 ), .IN6(n14386), .Q(n9457) );
  OR2X1 U1613 ( .IN1(n9459), .IN2(n9460), .Q(n9458) );
  AO221X1 U1614 ( .IN1(\U50/DATA1_10 ), .IN2(n14385), .IN3(
        p___constant_11x11xf32_10_1[10]), .IN4(n14373), .IN5(n9461), .Q(n9460)
         );
  AO22X1 U1615 ( .IN1(\U25/DATA1_10 ), .IN2(n14254), .IN3(
        p___constant_11x11xf32_10_0[10]), .IN4(n14360), .Q(n9461) );
  AO221X1 U1616 ( .IN1(\U30/DATA1_10 ), .IN2(n14354), .IN3(\U45/DATA1_10 ), 
        .IN4(n14343), .IN5(n9462), .Q(n9459) );
  AO22X1 U1617 ( .IN1(\U35/DATA1_10 ), .IN2(n14333), .IN3(\U40/DATA1_10 ), 
        .IN4(n14322), .Q(n9462) );
  AO221X1 U1618 ( .IN1(n14235), .IN2(n13967), .IN3(\U10/DATA1_9 ), .IN4(n14198), .IN5(n9464), .Q(n13139) );
  AO222X1 U1619 ( .IN1(p___constant_11x11xf32_10_9[9]), .IN2(n14407), .IN3(
        n14397), .IN4(n9465), .IN5(\U20/DATA1_9 ), .IN6(n14386), .Q(n9464) );
  OR2X1 U1620 ( .IN1(n9466), .IN2(n9467), .Q(n9465) );
  AO221X1 U1621 ( .IN1(\U50/DATA1_9 ), .IN2(n14385), .IN3(
        p___constant_11x11xf32_10_1[9]), .IN4(n14373), .IN5(n9468), .Q(n9467)
         );
  AO22X1 U1622 ( .IN1(\U25/DATA1_9 ), .IN2(n14256), .IN3(
        p___constant_11x11xf32_10_0[9]), .IN4(n14360), .Q(n9468) );
  AO221X1 U1623 ( .IN1(\U30/DATA1_9 ), .IN2(n14354), .IN3(\U45/DATA1_9 ), 
        .IN4(n14343), .IN5(n9469), .Q(n9466) );
  AO22X1 U1624 ( .IN1(\U35/DATA1_9 ), .IN2(n14333), .IN3(\U40/DATA1_9 ), .IN4(
        n14322), .Q(n9469) );
  AO221X1 U1626 ( .IN1(n14235), .IN2(\fmul_0_0_0_0_10/add_2_root_add_321/B[4] ), .IN3(p___constant_11x11xf32_10_10[8]), .IN4(n14200), .IN5(n9470), .Q(n13140)
         );
  AO222X1 U1627 ( .IN1(p___constant_11x11xf32_10_9[8]), .IN2(n14407), .IN3(
        n14397), .IN4(n9471), .IN5(\U20/DATA1_8 ), .IN6(n14386), .Q(n9470) );
  OR2X1 U1628 ( .IN1(n9472), .IN2(n9473), .Q(n9471) );
  AO221X1 U1629 ( .IN1(\U50/DATA1_8 ), .IN2(n14385), .IN3(
        p___constant_11x11xf32_10_1[8]), .IN4(n14373), .IN5(n9474), .Q(n9473)
         );
  AO22X1 U1630 ( .IN1(\U25/DATA1_8 ), .IN2(n14192), .IN3(
        p___constant_11x11xf32_10_0[8]), .IN4(n14360), .Q(n9474) );
  AO221X1 U1631 ( .IN1(p___constant_11x11xf32_10_6[8]), .IN2(n14354), .IN3(
        \U45/DATA1_8 ), .IN4(n14343), .IN5(n9475), .Q(n9472) );
  AO22X1 U1632 ( .IN1(\U35/DATA1_8 ), .IN2(n14333), .IN3(\U40/DATA1_8 ), .IN4(
        n14322), .Q(n9475) );
  AO221X1 U1633 ( .IN1(n14235), .IN2(\fmul_0_0_0_0_10/add_2_root_add_321/B[3] ), .IN3(p___constant_11x11xf32_10_10[7]), .IN4(n14199), .IN5(n9476), .Q(n13141)
         );
  AO222X1 U1634 ( .IN1(p___constant_11x11xf32_10_9[7]), .IN2(n14407), .IN3(
        n14397), .IN4(n9477), .IN5(\U20/DATA1_7 ), .IN6(n14386), .Q(n9476) );
  OR2X1 U1635 ( .IN1(n9478), .IN2(n9479), .Q(n9477) );
  AO221X1 U1636 ( .IN1(\U50/DATA1_7 ), .IN2(n14385), .IN3(
        p___constant_11x11xf32_10_1[7]), .IN4(n14373), .IN5(n9480), .Q(n9479)
         );
  AO22X1 U1637 ( .IN1(\U25/DATA1_7 ), .IN2(n14914), .IN3(
        p___constant_11x11xf32_10_0[7]), .IN4(n14360), .Q(n9480) );
  AO221X1 U1638 ( .IN1(p___constant_11x11xf32_10_6[7]), .IN2(n14354), .IN3(
        \U45/DATA1_7 ), .IN4(n14343), .IN5(n9481), .Q(n9478) );
  AO22X1 U1639 ( .IN1(\U35/DATA1_7 ), .IN2(n14333), .IN3(\U40/DATA1_7 ), .IN4(
        n14322), .Q(n9481) );
  AO221X1 U1640 ( .IN1(n14235), .IN2(\fmul_0_0_0_0_10/add_2_root_add_321/B[2] ), .IN3(p___constant_11x11xf32_10_10[6]), .IN4(n14194), .IN5(n9482), .Q(n13142)
         );
  AO222X1 U1641 ( .IN1(p___constant_11x11xf32_10_9[6]), .IN2(n14407), .IN3(
        n14397), .IN4(n9483), .IN5(\U20/DATA1_6 ), .IN6(n14386), .Q(n9482) );
  OR2X1 U1642 ( .IN1(n9484), .IN2(n9485), .Q(n9483) );
  AO221X1 U1643 ( .IN1(\U50/DATA1_6 ), .IN2(n14385), .IN3(
        p___constant_11x11xf32_10_1[6]), .IN4(n14373), .IN5(n9486), .Q(n9485)
         );
  AO22X1 U1644 ( .IN1(\U25/DATA1_6 ), .IN2(n14257), .IN3(
        p___constant_11x11xf32_10_0[6]), .IN4(n14360), .Q(n9486) );
  AO221X1 U1645 ( .IN1(p___constant_11x11xf32_10_6[6]), .IN2(n14354), .IN3(
        \U45/DATA1_6 ), .IN4(n14343), .IN5(n9487), .Q(n9484) );
  AO22X1 U1646 ( .IN1(\U35/DATA1_6 ), .IN2(n14333), .IN3(\U40/DATA1_6 ), .IN4(
        n14322), .Q(n9487) );
  AO221X1 U1647 ( .IN1(n14235), .IN2(\fmul_0_0_0_0_10/add_2_root_add_321/B[1] ), .IN3(p___constant_11x11xf32_10_10[5]), .IN4(n14195), .IN5(n9488), .Q(n13143)
         );
  AO222X1 U1648 ( .IN1(p___constant_11x11xf32_10_9[5]), .IN2(n14407), .IN3(
        n14397), .IN4(n9489), .IN5(p___constant_11x11xf32_10_8[5]), .IN6(
        n14386), .Q(n9488) );
  OR2X1 U1649 ( .IN1(n9490), .IN2(n9491), .Q(n9489) );
  AO221X1 U1650 ( .IN1(\U50/DATA1_5 ), .IN2(n14385), .IN3(
        p___constant_11x11xf32_10_1[5]), .IN4(n14373), .IN5(n9492), .Q(n9491)
         );
  AO22X1 U1651 ( .IN1(\U25/DATA1_5 ), .IN2(n14257), .IN3(
        p___constant_11x11xf32_10_0[5]), .IN4(n14360), .Q(n9492) );
  AO221X1 U1652 ( .IN1(p___constant_11x11xf32_10_6[5]), .IN2(n14354), .IN3(
        \U45/DATA1_5 ), .IN4(n14343), .IN5(n9493), .Q(n9490) );
  AO22X1 U1653 ( .IN1(\U35/DATA1_5 ), .IN2(n14333), .IN3(\U40/DATA1_5 ), .IN4(
        n14322), .Q(n9493) );
  AO221X1 U1654 ( .IN1(n14235), .IN2(\fmul_0_0_0_0_10/add_2_root_add_321/B[0] ), .IN3(p___constant_11x11xf32_10_10[4]), .IN4(n14197), .IN5(n9494), .Q(n13144)
         );
  AO222X1 U1655 ( .IN1(p___constant_11x11xf32_10_9[4]), .IN2(n14407), .IN3(
        n14397), .IN4(n9495), .IN5(p___constant_11x11xf32_10_8[4]), .IN6(
        n14386), .Q(n9494) );
  OR2X1 U1656 ( .IN1(n9496), .IN2(n9497), .Q(n9495) );
  AO221X1 U1657 ( .IN1(\U50/DATA1_4 ), .IN2(n14385), .IN3(
        p___constant_11x11xf32_10_1[4]), .IN4(n14373), .IN5(n9498), .Q(n9497)
         );
  AO22X1 U1658 ( .IN1(\U25/DATA1_4 ), .IN2(n14256), .IN3(
        p___constant_11x11xf32_10_0[4]), .IN4(n14360), .Q(n9498) );
  AO221X1 U1659 ( .IN1(p___constant_11x11xf32_10_6[4]), .IN2(n14354), .IN3(
        p___constant_11x11xf32_10_3[4]), .IN4(n14343), .IN5(n9499), .Q(n9496)
         );
  AO22X1 U1660 ( .IN1(\U35/DATA1_4 ), .IN2(n14333), .IN3(\U40/DATA1_4 ), .IN4(
        n14322), .Q(n9499) );
  AO221X1 U1661 ( .IN1(n14235), .IN2(n13499), .IN3(
        p___constant_11x11xf32_10_10[3]), .IN4(n14196), .IN5(n9501), .Q(n13145) );
  AO222X1 U1662 ( .IN1(p___constant_11x11xf32_10_9[3]), .IN2(n14407), .IN3(
        n14397), .IN4(n9502), .IN5(p___constant_11x11xf32_10_8[3]), .IN6(
        n14386), .Q(n9501) );
  OR2X1 U1663 ( .IN1(n9503), .IN2(n9504), .Q(n9502) );
  AO221X1 U1664 ( .IN1(p___constant_11x11xf32_10_2[3]), .IN2(n14385), .IN3(
        p___constant_11x11xf32_10_1[3]), .IN4(n14373), .IN5(n9505), .Q(n9504)
         );
  AO22X1 U1665 ( .IN1(\U25/DATA1_3 ), .IN2(n14189), .IN3(
        p___constant_11x11xf32_10_0[3]), .IN4(n14360), .Q(n9505) );
  AO221X1 U1666 ( .IN1(p___constant_11x11xf32_10_6[3]), .IN2(n14354), .IN3(
        p___constant_11x11xf32_10_3[3]), .IN4(n14343), .IN5(n9506), .Q(n9503)
         );
  AO22X1 U1667 ( .IN1(p___constant_11x11xf32_10_5[3]), .IN2(n14333), .IN3(
        \U40/DATA1_3 ), .IN4(n14322), .Q(n9506) );
  AO221X1 U1668 ( .IN1(n14235), .IN2(n13617), .IN3(
        p___constant_11x11xf32_10_10[2]), .IN4(n14198), .IN5(n9508), .Q(n13146) );
  AO222X1 U1669 ( .IN1(p___constant_11x11xf32_10_9[2]), .IN2(n14407), .IN3(
        n14397), .IN4(n9509), .IN5(p___constant_11x11xf32_10_8[2]), .IN6(
        n14386), .Q(n9508) );
  OR2X1 U1670 ( .IN1(n9510), .IN2(n9511), .Q(n9509) );
  AO221X1 U1671 ( .IN1(p___constant_11x11xf32_10_2[2]), .IN2(n14385), .IN3(
        p___constant_11x11xf32_10_1[2]), .IN4(n14373), .IN5(n9512), .Q(n9511)
         );
  AO22X1 U1672 ( .IN1(\U25/DATA1_2 ), .IN2(n14254), .IN3(
        p___constant_11x11xf32_10_0[2]), .IN4(n14360), .Q(n9512) );
  AO221X1 U1673 ( .IN1(p___constant_11x11xf32_10_6[2]), .IN2(n14354), .IN3(
        p___constant_11x11xf32_10_3[2]), .IN4(n14343), .IN5(n9513), .Q(n9510)
         );
  AO22X1 U1674 ( .IN1(p___constant_11x11xf32_10_5[2]), .IN2(n14333), .IN3(
        \U40/DATA1_2 ), .IN4(n14322), .Q(n9513) );
  AO221X1 U1675 ( .IN1(n14235), .IN2(n13620), .IN3(
        p___constant_11x11xf32_10_10[1]), .IN4(n14200), .IN5(n9515), .Q(n13147) );
  AO222X1 U1676 ( .IN1(p___constant_11x11xf32_10_9[1]), .IN2(n14407), .IN3(
        n14397), .IN4(n9516), .IN5(p___constant_11x11xf32_10_8[1]), .IN6(
        n14386), .Q(n9515) );
  OR2X1 U1677 ( .IN1(n9517), .IN2(n9518), .Q(n9516) );
  AO221X1 U1678 ( .IN1(p___constant_11x11xf32_10_2[1]), .IN2(n14385), .IN3(
        p___constant_11x11xf32_10_1[1]), .IN4(n14373), .IN5(n9519), .Q(n9518)
         );
  AO22X1 U1679 ( .IN1(\U25/DATA1_1 ), .IN2(n14186), .IN3(
        p___constant_11x11xf32_10_0[1]), .IN4(n14359), .Q(n9519) );
  AO221X1 U1680 ( .IN1(p___constant_11x11xf32_10_6[1]), .IN2(n14354), .IN3(
        p___constant_11x11xf32_10_3[1]), .IN4(n14343), .IN5(n9520), .Q(n9517)
         );
  AO22X1 U1681 ( .IN1(p___constant_11x11xf32_10_5[1]), .IN2(n14333), .IN3(
        \U40/DATA1_1 ), .IN4(n14322), .Q(n9520) );
  AO221X1 U1682 ( .IN1(n14236), .IN2(n13618), .IN3(
        p___constant_11x11xf32_10_10[0]), .IN4(n14199), .IN5(n9522), .Q(n13148) );
  AO222X1 U1683 ( .IN1(p___constant_11x11xf32_10_9[0]), .IN2(n14407), .IN3(
        n14397), .IN4(n9523), .IN5(p___constant_11x11xf32_10_8[0]), .IN6(
        n14386), .Q(n9522) );
  OR2X1 U1684 ( .IN1(n9524), .IN2(n9525), .Q(n9523) );
  AO221X1 U1685 ( .IN1(p___constant_11x11xf32_10_2[0]), .IN2(n14385), .IN3(
        p___constant_11x11xf32_10_1[0]), .IN4(n14373), .IN5(n9526), .Q(n9525)
         );
  AO22X1 U1686 ( .IN1(p___constant_11x11xf32_10_7[0]), .IN2(n14190), .IN3(
        p___constant_11x11xf32_10_0[0]), .IN4(n14359), .Q(n9526) );
  AO221X1 U1687 ( .IN1(p___constant_11x11xf32_10_6[0]), .IN2(n14354), .IN3(
        p___constant_11x11xf32_10_3[0]), .IN4(n14343), .IN5(n9527), .Q(n9524)
         );
  AO22X1 U1688 ( .IN1(p___constant_11x11xf32_10_5[0]), .IN2(n14333), .IN3(
        p___constant_11x11xf32_10_4[0]), .IN4(n14322), .Q(n9527) );
  AO21X1 U1689 ( .IN1(n14238), .IN2(n13765), .IN3(n9529), .Q(n13149) );
  AO21X1 U1690 ( .IN1(n14239), .IN2(n13897), .IN3(n9531), .Q(n13150) );
  AO21X1 U1691 ( .IN1(n14238), .IN2(n14077), .IN3(n9533), .Q(n13151) );
  AO21X1 U1693 ( .IN1(n14238), .IN2(\fmul_0_0_0_0_10/add_2_root_add_321/A[4] ), 
        .IN3(n9534), .Q(n13152) );
  AO21X1 U1694 ( .IN1(n14239), .IN2(\fmul_0_0_0_0_10/add_2_root_add_321/A[3] ), 
        .IN3(n9535), .Q(n13153) );
  AO21X1 U1695 ( .IN1(n14238), .IN2(\fmul_0_0_0_0_10/add_2_root_add_321/A[2] ), 
        .IN3(n9536), .Q(n13154) );
  AO21X1 U1696 ( .IN1(n14238), .IN2(\fmul_0_0_0_0_10/add_2_root_add_321/A[1] ), 
        .IN3(n9537), .Q(n13155) );
  AO21X1 U1697 ( .IN1(n14239), .IN2(\fmul_0_0_0_0_10/add_2_root_add_321/A[0] ), 
        .IN3(n9538), .Q(n13156) );
  AO21X1 U1698 ( .IN1(n14239), .IN2(n13468), .IN3(n9540), .Q(n13157) );
  AO21X1 U1699 ( .IN1(n14239), .IN2(n13619), .IN3(n9542), .Q(n13158) );
  AO21X1 U1700 ( .IN1(n14239), .IN2(n13629), .IN3(n9544), .Q(n13159) );
  AO221X1 U1702 ( .IN1(n14236), .IN2(n13907), .IN3(\U63/DATA1_11 ), .IN4(
        n14194), .IN5(n9546), .Q(n13161) );
  AO222X1 U1703 ( .IN1(\U68/DATA1_11 ), .IN2(n14407), .IN3(n14398), .IN4(n9547), .IN5(\U73/DATA1_11 ), .IN6(n14387), .Q(n9546) );
  OR2X1 U1704 ( .IN1(n9548), .IN2(n9549), .Q(n9547) );
  AO221X1 U1705 ( .IN1(\U103/DATA1_11 ), .IN2(n14384), .IN3(\U108/DATA1_11 ), 
        .IN4(n14372), .IN5(n9550), .Q(n9549) );
  AO22X1 U1706 ( .IN1(\U78/DATA1_11 ), .IN2(n14254), .IN3(\U108/DATA2_11 ), 
        .IN4(n14359), .Q(n9550) );
  AO221X1 U1707 ( .IN1(\U83/DATA1_11 ), .IN2(n14353), .IN3(\U98/DATA1_11 ), 
        .IN4(n14342), .IN5(n9551), .Q(n9548) );
  AO22X1 U1708 ( .IN1(\U88/DATA1_11 ), .IN2(n14332), .IN3(\U93/DATA1_11 ), 
        .IN4(n14321), .Q(n9551) );
  AO221X1 U1710 ( .IN1(n14236), .IN2(n13606), .IN3(
        p___constant_11x11xf32_9_10[10]), .IN4(n14195), .IN5(n9553), .Q(n13162) );
  AO222X1 U1711 ( .IN1(\U68/DATA1_10 ), .IN2(n14407), .IN3(n14398), .IN4(n9554), .IN5(\U73/DATA1_10 ), .IN6(n14387), .Q(n9553) );
  OR2X1 U1712 ( .IN1(n9555), .IN2(n9556), .Q(n9554) );
  AO221X1 U1713 ( .IN1(\U103/DATA1_10 ), .IN2(n14384), .IN3(\U108/DATA1_10 ), 
        .IN4(n14372), .IN5(n9557), .Q(n9556) );
  AO22X1 U1714 ( .IN1(\U78/DATA1_10 ), .IN2(n14254), .IN3(\U108/DATA2_10 ), 
        .IN4(n14359), .Q(n9557) );
  AO221X1 U1715 ( .IN1(\U83/DATA1_10 ), .IN2(n14353), .IN3(\U98/DATA1_10 ), 
        .IN4(n14342), .IN5(n9558), .Q(n9555) );
  AO22X1 U1716 ( .IN1(\U88/DATA1_10 ), .IN2(n14332), .IN3(\U93/DATA1_10 ), 
        .IN4(n14321), .Q(n9558) );
  AO221X1 U1717 ( .IN1(n14237), .IN2(n13966), .IN3(
        p___constant_11x11xf32_9_10[9]), .IN4(n14197), .IN5(n9560), .Q(n13163)
         );
  AO222X1 U1718 ( .IN1(\U68/DATA1_9 ), .IN2(n14407), .IN3(n14398), .IN4(n9561), 
        .IN5(\U73/DATA1_9 ), .IN6(n14387), .Q(n9560) );
  OR2X1 U1719 ( .IN1(n9562), .IN2(n9563), .Q(n9561) );
  AO221X1 U1720 ( .IN1(\U103/DATA1_9 ), .IN2(n14384), .IN3(\U108/DATA1_9 ), 
        .IN4(n14372), .IN5(n9564), .Q(n9563) );
  AO22X1 U1721 ( .IN1(\U78/DATA1_9 ), .IN2(n14254), .IN3(\U108/DATA2_9 ), 
        .IN4(n14359), .Q(n9564) );
  AO221X1 U1722 ( .IN1(\U83/DATA1_9 ), .IN2(n14353), .IN3(\U98/DATA1_9 ), 
        .IN4(n14342), .IN5(n9565), .Q(n9562) );
  AO22X1 U1723 ( .IN1(\U88/DATA1_9 ), .IN2(n14332), .IN3(\U93/DATA1_9 ), .IN4(
        n14321), .Q(n9565) );
  AO221X1 U1725 ( .IN1(n5302), .IN2(n14247), .IN3(
        p___constant_11x11xf32_9_10[8]), .IN4(n14196), .IN5(n9566), .Q(n13164)
         );
  AO222X1 U1726 ( .IN1(\U68/DATA1_8 ), .IN2(n14407), .IN3(n14398), .IN4(n9567), 
        .IN5(\U73/DATA1_8 ), .IN6(n14387), .Q(n9566) );
  OR2X1 U1727 ( .IN1(n9568), .IN2(n9569), .Q(n9567) );
  AO221X1 U1728 ( .IN1(\U103/DATA1_8 ), .IN2(n14384), .IN3(\U108/DATA1_8 ), 
        .IN4(n14372), .IN5(n9570), .Q(n9569) );
  AO22X1 U1729 ( .IN1(p___constant_11x11xf32_9_7[8]), .IN2(n14186), .IN3(
        \U108/DATA2_8 ), .IN4(n14359), .Q(n9570) );
  AO221X1 U1730 ( .IN1(\U83/DATA1_8 ), .IN2(n14353), .IN3(\U98/DATA1_8 ), 
        .IN4(n14342), .IN5(n9571), .Q(n9568) );
  AO22X1 U1731 ( .IN1(\U88/DATA1_8 ), .IN2(n14332), .IN3(\U93/DATA1_8 ), .IN4(
        n14321), .Q(n9571) );
  AO221X1 U1732 ( .IN1(n5301), .IN2(n14247), .IN3(
        p___constant_11x11xf32_9_10[7]), .IN4(n14198), .IN5(n9572), .Q(n13165)
         );
  AO222X1 U1733 ( .IN1(\U68/DATA1_7 ), .IN2(n14408), .IN3(n14398), .IN4(n9573), 
        .IN5(\U73/DATA1_7 ), .IN6(n14387), .Q(n9572) );
  OR2X1 U1734 ( .IN1(n9574), .IN2(n9575), .Q(n9573) );
  AO221X1 U1735 ( .IN1(\U103/DATA1_7 ), .IN2(n14384), .IN3(\U108/DATA1_7 ), 
        .IN4(n14372), .IN5(n9576), .Q(n9575) );
  AO22X1 U1736 ( .IN1(p___constant_11x11xf32_9_7[7]), .IN2(n14190), .IN3(
        \U108/DATA2_7 ), .IN4(n14359), .Q(n9576) );
  AO221X1 U1737 ( .IN1(\U83/DATA1_7 ), .IN2(n14353), .IN3(\U98/DATA1_7 ), 
        .IN4(n14342), .IN5(n9577), .Q(n9574) );
  AO22X1 U1738 ( .IN1(\U88/DATA1_7 ), .IN2(n14332), .IN3(\U93/DATA1_7 ), .IN4(
        n14321), .Q(n9577) );
  AO221X1 U1739 ( .IN1(n5300), .IN2(n14247), .IN3(
        p___constant_11x11xf32_9_10[6]), .IN4(n14200), .IN5(n9578), .Q(n13166)
         );
  AO222X1 U1740 ( .IN1(\U68/DATA1_6 ), .IN2(n14408), .IN3(n14398), .IN4(n9579), 
        .IN5(\U73/DATA1_6 ), .IN6(n14387), .Q(n9578) );
  OR2X1 U1741 ( .IN1(n9580), .IN2(n9581), .Q(n9579) );
  AO221X1 U1742 ( .IN1(\U103/DATA1_6 ), .IN2(n14384), .IN3(\U108/DATA1_6 ), 
        .IN4(n14372), .IN5(n9582), .Q(n9581) );
  AO22X1 U1743 ( .IN1(p___constant_11x11xf32_9_7[6]), .IN2(n14193), .IN3(
        \U108/DATA2_6 ), .IN4(n14359), .Q(n9582) );
  AO221X1 U1744 ( .IN1(\U83/DATA1_6 ), .IN2(n14353), .IN3(\U98/DATA1_6 ), 
        .IN4(n14342), .IN5(n9583), .Q(n9580) );
  AO22X1 U1745 ( .IN1(\U88/DATA1_6 ), .IN2(n14332), .IN3(\U93/DATA1_6 ), .IN4(
        n14321), .Q(n9583) );
  AO221X1 U1746 ( .IN1(n5299), .IN2(n14247), .IN3(
        p___constant_11x11xf32_9_10[5]), .IN4(n14199), .IN5(n9584), .Q(n13167)
         );
  AO222X1 U1747 ( .IN1(p___constant_11x11xf32_9_9[5]), .IN2(n14408), .IN3(
        n14398), .IN4(n9585), .IN5(\U73/DATA1_5 ), .IN6(n14387), .Q(n9584) );
  OR2X1 U1748 ( .IN1(n9586), .IN2(n9587), .Q(n9585) );
  AO221X1 U1749 ( .IN1(\U103/DATA1_5 ), .IN2(n14384), .IN3(\U108/DATA1_5 ), 
        .IN4(n14372), .IN5(n9588), .Q(n9587) );
  AO22X1 U1750 ( .IN1(p___constant_11x11xf32_9_7[5]), .IN2(n14257), .IN3(
        \U108/DATA2_5 ), .IN4(n14359), .Q(n9588) );
  AO221X1 U1751 ( .IN1(\U83/DATA1_5 ), .IN2(n14353), .IN3(\U98/DATA1_5 ), 
        .IN4(n14342), .IN5(n9589), .Q(n9586) );
  AO22X1 U1752 ( .IN1(\U88/DATA1_5 ), .IN2(n14332), .IN3(\U93/DATA1_5 ), .IN4(
        n14321), .Q(n9589) );
  AO221X1 U1753 ( .IN1(n5298), .IN2(n14248), .IN3(
        p___constant_11x11xf32_9_10[4]), .IN4(n14194), .IN5(n9590), .Q(n13168)
         );
  AO222X1 U1754 ( .IN1(p___constant_11x11xf32_9_9[4]), .IN2(n14408), .IN3(
        n14398), .IN4(n9591), .IN5(\U73/DATA1_4 ), .IN6(n14387), .Q(n9590) );
  OR2X1 U1755 ( .IN1(n9592), .IN2(n9593), .Q(n9591) );
  AO221X1 U1756 ( .IN1(\U103/DATA1_4 ), .IN2(n14384), .IN3(\U108/DATA1_4 ), 
        .IN4(n14372), .IN5(n9594), .Q(n9593) );
  AO22X1 U1757 ( .IN1(p___constant_11x11xf32_9_7[4]), .IN2(n14189), .IN3(
        \U108/DATA2_4 ), .IN4(n14359), .Q(n9594) );
  AO221X1 U1758 ( .IN1(\U83/DATA1_4 ), .IN2(n14353), .IN3(\U98/DATA1_4 ), 
        .IN4(n14342), .IN5(n9595), .Q(n9592) );
  AO22X1 U1759 ( .IN1(\U88/DATA1_4 ), .IN2(n14332), .IN3(
        p___constant_11x11xf32_9_4[4]), .IN4(n14321), .Q(n9595) );
  AO221X1 U1760 ( .IN1(n5297), .IN2(n14248), .IN3(
        p___constant_11x11xf32_9_10[3]), .IN4(n14195), .IN5(n9596), .Q(n13169)
         );
  AO222X1 U1761 ( .IN1(p___constant_11x11xf32_9_9[3]), .IN2(n14408), .IN3(
        n14398), .IN4(n9597), .IN5(\U73/DATA1_3 ), .IN6(n14387), .Q(n9596) );
  OR2X1 U1762 ( .IN1(n9598), .IN2(n9599), .Q(n9597) );
  AO221X1 U1763 ( .IN1(\U103/DATA1_3 ), .IN2(n14384), .IN3(\U108/DATA1_3 ), 
        .IN4(n14372), .IN5(n9600), .Q(n9599) );
  AO22X1 U1764 ( .IN1(p___constant_11x11xf32_9_7[3]), .IN2(n14191), .IN3(
        \U108/DATA2_3 ), .IN4(n14359), .Q(n9600) );
  AO221X1 U1765 ( .IN1(p___constant_11x11xf32_9_6[3]), .IN2(n14353), .IN3(
        \U98/DATA1_3 ), .IN4(n14342), .IN5(n9601), .Q(n9598) );
  AO22X1 U1766 ( .IN1(\U88/DATA1_3 ), .IN2(n14332), .IN3(
        p___constant_11x11xf32_9_4[3]), .IN4(n14321), .Q(n9601) );
  AO221X1 U1767 ( .IN1(n5296), .IN2(n14248), .IN3(
        p___constant_11x11xf32_9_10[2]), .IN4(n14197), .IN5(n9602), .Q(n13170)
         );
  AO222X1 U1768 ( .IN1(p___constant_11x11xf32_9_9[2]), .IN2(n14408), .IN3(
        n14398), .IN4(n9603), .IN5(\U73/DATA1_2 ), .IN6(n14387), .Q(n9602) );
  OR2X1 U1769 ( .IN1(n9604), .IN2(n9605), .Q(n9603) );
  AO221X1 U1770 ( .IN1(\U103/DATA1_2 ), .IN2(n14384), .IN3(\U108/DATA1_2 ), 
        .IN4(n14372), .IN5(n9606), .Q(n9605) );
  AO22X1 U1771 ( .IN1(p___constant_11x11xf32_9_7[2]), .IN2(n14914), .IN3(
        \U108/DATA2_2 ), .IN4(n14359), .Q(n9606) );
  AO221X1 U1772 ( .IN1(p___constant_11x11xf32_9_6[2]), .IN2(n14353), .IN3(
        \U98/DATA1_2 ), .IN4(n14342), .IN5(n9607), .Q(n9604) );
  AO22X1 U1773 ( .IN1(\U88/DATA1_2 ), .IN2(n14332), .IN3(
        p___constant_11x11xf32_9_4[2]), .IN4(n14321), .Q(n9607) );
  AO221X1 U1774 ( .IN1(n5295), .IN2(n14248), .IN3(
        p___constant_11x11xf32_9_10[1]), .IN4(n14196), .IN5(n9608), .Q(n13171)
         );
  AO222X1 U1775 ( .IN1(p___constant_11x11xf32_9_9[1]), .IN2(n14408), .IN3(
        n14398), .IN4(n9609), .IN5(\U73/DATA1_1 ), .IN6(n14387), .Q(n9608) );
  OR2X1 U1776 ( .IN1(n9610), .IN2(n9611), .Q(n9609) );
  AO221X1 U1777 ( .IN1(\U103/DATA1_1 ), .IN2(n14384), .IN3(\U108/DATA1_1 ), 
        .IN4(n14372), .IN5(n9612), .Q(n9611) );
  AO22X1 U1778 ( .IN1(p___constant_11x11xf32_9_7[1]), .IN2(n14186), .IN3(
        \U108/DATA2_1 ), .IN4(n14359), .Q(n9612) );
  AO221X1 U1779 ( .IN1(p___constant_11x11xf32_9_6[1]), .IN2(n14353), .IN3(
        \U98/DATA1_1 ), .IN4(n14342), .IN5(n9613), .Q(n9610) );
  AO22X1 U1780 ( .IN1(\U88/DATA1_1 ), .IN2(n14332), .IN3(
        p___constant_11x11xf32_9_4[1]), .IN4(n14321), .Q(n9613) );
  AO221X1 U1781 ( .IN1(n5294), .IN2(n14248), .IN3(
        p___constant_11x11xf32_9_10[0]), .IN4(n14198), .IN5(n9614), .Q(n13172)
         );
  AO222X1 U1782 ( .IN1(p___constant_11x11xf32_9_9[0]), .IN2(n14408), .IN3(
        n14398), .IN4(n9615), .IN5(p___constant_11x11xf32_9_8[0]), .IN6(n14387), .Q(n9614) );
  OR2X1 U1783 ( .IN1(n9616), .IN2(n9617), .Q(n9615) );
  AO221X1 U1784 ( .IN1(\U103/DATA1_0 ), .IN2(n14384), .IN3(\U108/DATA1_0 ), 
        .IN4(n14372), .IN5(n9618), .Q(n9617) );
  AO22X1 U1785 ( .IN1(p___constant_11x11xf32_9_7[0]), .IN2(n14914), .IN3(
        \U108/DATA2_0 ), .IN4(n14359), .Q(n9618) );
  AO221X1 U1786 ( .IN1(p___constant_11x11xf32_9_6[0]), .IN2(n14353), .IN3(
        \U98/DATA1_0 ), .IN4(n14342), .IN5(n9619), .Q(n9616) );
  AO22X1 U1787 ( .IN1(p___constant_11x11xf32_9_5[0]), .IN2(n14332), .IN3(
        p___constant_11x11xf32_9_4[0]), .IN4(n14321), .Q(n9619) );
  AO21X1 U1788 ( .IN1(n14239), .IN2(n13764), .IN3(n9529), .Q(n13173) );
  AO21X1 U1789 ( .IN1(n14238), .IN2(n13896), .IN3(n9531), .Q(n13174) );
  AO21X1 U1790 ( .IN1(n14240), .IN2(n14076), .IN3(n9533), .Q(n13175) );
  AO21X1 U1792 ( .IN1(n5314), .IN2(n14244), .IN3(n9534), .Q(n13176) );
  AO21X1 U1793 ( .IN1(n5313), .IN2(n14244), .IN3(n9535), .Q(n13177) );
  AO21X1 U1794 ( .IN1(n5312), .IN2(n14244), .IN3(n9536), .Q(n13178) );
  AO21X1 U1795 ( .IN1(n5311), .IN2(n14244), .IN3(n9537), .Q(n13179) );
  AO21X1 U1796 ( .IN1(n5310), .IN2(n14244), .IN3(n9538), .Q(n13180) );
  AO21X1 U1797 ( .IN1(n5309), .IN2(n14244), .IN3(n9540), .Q(n13181) );
  AO21X1 U1798 ( .IN1(n5308), .IN2(n14244), .IN3(n9542), .Q(n13182) );
  AO21X1 U1799 ( .IN1(n5307), .IN2(n14243), .IN3(n9544), .Q(n13183) );
  AO221X1 U1801 ( .IN1(n14235), .IN2(n13906), .IN3(\U125/DATA1_11 ), .IN4(
        n14200), .IN5(n9624), .Q(n13185) );
  AO222X1 U1802 ( .IN1(\U130/DATA1_11 ), .IN2(n14408), .IN3(n14399), .IN4(
        n9625), .IN5(\U135/DATA1_11 ), .IN6(n14388), .Q(n9624) );
  OR2X1 U1803 ( .IN1(n9626), .IN2(n9627), .Q(n9625) );
  AO221X1 U1804 ( .IN1(\U165/DATA1_11 ), .IN2(n14383), .IN3(\U170/DATA1_11 ), 
        .IN4(n14371), .IN5(n9628), .Q(n9627) );
  AO22X1 U1805 ( .IN1(\U140/DATA1_11 ), .IN2(n14254), .IN3(\U170/DATA2_11 ), 
        .IN4(n14359), .Q(n9628) );
  AO221X1 U1806 ( .IN1(\U145/DATA1_11 ), .IN2(n14352), .IN3(\U160/DATA1_11 ), 
        .IN4(n14341), .IN5(n9629), .Q(n9626) );
  AO22X1 U1807 ( .IN1(\U150/DATA1_11 ), .IN2(n14331), .IN3(\U155/DATA1_11 ), 
        .IN4(n14321), .Q(n9629) );
  AO221X1 U1809 ( .IN1(n14236), .IN2(n13605), .IN3(\U125/DATA1_10 ), .IN4(
        n14200), .IN5(n9631), .Q(n13186) );
  AO222X1 U1810 ( .IN1(\U130/DATA1_10 ), .IN2(n14408), .IN3(n14399), .IN4(
        n9632), .IN5(\U135/DATA1_10 ), .IN6(n14388), .Q(n9631) );
  OR2X1 U1811 ( .IN1(n9633), .IN2(n9634), .Q(n9632) );
  AO221X1 U1812 ( .IN1(\U165/DATA1_10 ), .IN2(n14383), .IN3(\U170/DATA1_10 ), 
        .IN4(n14371), .IN5(n9635), .Q(n9634) );
  AO22X1 U1813 ( .IN1(\U140/DATA1_10 ), .IN2(n14193), .IN3(\U170/DATA2_10 ), 
        .IN4(n14358), .Q(n9635) );
  AO221X1 U1814 ( .IN1(\U145/DATA1_10 ), .IN2(n14352), .IN3(\U160/DATA1_10 ), 
        .IN4(n14341), .IN5(n9636), .Q(n9633) );
  AO22X1 U1815 ( .IN1(\U150/DATA1_10 ), .IN2(n14331), .IN3(\U155/DATA1_10 ), 
        .IN4(n14322), .Q(n9636) );
  AO221X1 U1816 ( .IN1(n14237), .IN2(n13965), .IN3(\U125/DATA1_9 ), .IN4(
        n14200), .IN5(n9638), .Q(n13187) );
  AO222X1 U1817 ( .IN1(\U130/DATA1_9 ), .IN2(n14408), .IN3(n14399), .IN4(n9639), .IN5(\U135/DATA1_9 ), .IN6(n14388), .Q(n9638) );
  OR2X1 U1818 ( .IN1(n9640), .IN2(n9641), .Q(n9639) );
  AO221X1 U1819 ( .IN1(\U165/DATA1_9 ), .IN2(n14383), .IN3(\U170/DATA1_9 ), 
        .IN4(n14371), .IN5(n9642), .Q(n9641) );
  AO22X1 U1820 ( .IN1(\U140/DATA1_9 ), .IN2(n14257), .IN3(\U170/DATA2_9 ), 
        .IN4(n14358), .Q(n9642) );
  AO221X1 U1821 ( .IN1(\U145/DATA1_9 ), .IN2(n14352), .IN3(\U160/DATA1_9 ), 
        .IN4(n14341), .IN5(n9643), .Q(n9640) );
  AO22X1 U1822 ( .IN1(\U150/DATA1_9 ), .IN2(n14331), .IN3(\U155/DATA1_9 ), 
        .IN4(n14315), .Q(n9643) );
  AO221X1 U1824 ( .IN1(n5374), .IN2(n14249), .IN3(\U125/DATA1_8 ), .IN4(n14200), .IN5(n9644), .Q(n13188) );
  AO222X1 U1825 ( .IN1(\U130/DATA1_8 ), .IN2(n14408), .IN3(n14399), .IN4(n9645), .IN5(\U135/DATA1_8 ), .IN6(n14388), .Q(n9644) );
  OR2X1 U1826 ( .IN1(n9646), .IN2(n9647), .Q(n9645) );
  AO221X1 U1827 ( .IN1(\U165/DATA1_8 ), .IN2(n14383), .IN3(\U170/DATA1_8 ), 
        .IN4(n14371), .IN5(n9648), .Q(n9647) );
  AO22X1 U1828 ( .IN1(\U140/DATA1_8 ), .IN2(n14255), .IN3(\U170/DATA2_8 ), 
        .IN4(n14358), .Q(n9648) );
  AO221X1 U1829 ( .IN1(\U145/DATA1_8 ), .IN2(n14352), .IN3(\U160/DATA1_8 ), 
        .IN4(n14341), .IN5(n9649), .Q(n9646) );
  AO22X1 U1830 ( .IN1(\U150/DATA1_8 ), .IN2(n14331), .IN3(\U155/DATA1_8 ), 
        .IN4(n14315), .Q(n9649) );
  AO221X1 U1831 ( .IN1(n5373), .IN2(n14249), .IN3(\U125/DATA1_7 ), .IN4(n14200), .IN5(n9650), .Q(n13189) );
  AO222X1 U1832 ( .IN1(\U130/DATA1_7 ), .IN2(n14408), .IN3(n14399), .IN4(n9651), .IN5(\U135/DATA1_7 ), .IN6(n14388), .Q(n9650) );
  OR2X1 U1833 ( .IN1(n9652), .IN2(n9653), .Q(n9651) );
  AO221X1 U1834 ( .IN1(\U165/DATA1_7 ), .IN2(n14383), .IN3(\U170/DATA1_7 ), 
        .IN4(n14371), .IN5(n9654), .Q(n9653) );
  AO22X1 U1835 ( .IN1(\U140/DATA1_7 ), .IN2(n14191), .IN3(\U170/DATA2_7 ), 
        .IN4(n14358), .Q(n9654) );
  AO221X1 U1836 ( .IN1(\U145/DATA1_7 ), .IN2(n14352), .IN3(\U160/DATA1_7 ), 
        .IN4(n14341), .IN5(n9655), .Q(n9652) );
  AO22X1 U1837 ( .IN1(\U150/DATA1_7 ), .IN2(n14331), .IN3(\U155/DATA1_7 ), 
        .IN4(n14316), .Q(n9655) );
  AO221X1 U1838 ( .IN1(n5372), .IN2(n14249), .IN3(\U125/DATA1_6 ), .IN4(n14194), .IN5(n9656), .Q(n13190) );
  AO222X1 U1839 ( .IN1(\U130/DATA1_6 ), .IN2(n14408), .IN3(n14399), .IN4(n9657), .IN5(\U135/DATA1_6 ), .IN6(n14388), .Q(n9656) );
  OR2X1 U1840 ( .IN1(n9658), .IN2(n9659), .Q(n9657) );
  AO221X1 U1841 ( .IN1(\U165/DATA1_6 ), .IN2(n14383), .IN3(\U170/DATA1_6 ), 
        .IN4(n14371), .IN5(n9660), .Q(n9659) );
  AO22X1 U1842 ( .IN1(\U140/DATA1_6 ), .IN2(n14193), .IN3(\U170/DATA2_6 ), 
        .IN4(n14358), .Q(n9660) );
  AO221X1 U1843 ( .IN1(\U145/DATA1_6 ), .IN2(n14352), .IN3(\U160/DATA1_6 ), 
        .IN4(n14341), .IN5(n9661), .Q(n9658) );
  AO22X1 U1844 ( .IN1(\U150/DATA1_6 ), .IN2(n14331), .IN3(\U155/DATA1_6 ), 
        .IN4(n14320), .Q(n9661) );
  AO221X1 U1845 ( .IN1(n5371), .IN2(n14249), .IN3(\U125/DATA1_5 ), .IN4(n14194), .IN5(n9662), .Q(n13191) );
  AO222X1 U1846 ( .IN1(\U130/DATA1_5 ), .IN2(n14408), .IN3(n14399), .IN4(n9663), .IN5(\U135/DATA1_5 ), .IN6(n14388), .Q(n9662) );
  OR2X1 U1847 ( .IN1(n9664), .IN2(n9665), .Q(n9663) );
  AO221X1 U1848 ( .IN1(\U165/DATA1_5 ), .IN2(n14383), .IN3(\U170/DATA1_5 ), 
        .IN4(n14371), .IN5(n9666), .Q(n9665) );
  AO22X1 U1849 ( .IN1(\U140/DATA1_5 ), .IN2(n14257), .IN3(\U170/DATA2_5 ), 
        .IN4(n14358), .Q(n9666) );
  AO221X1 U1850 ( .IN1(\U145/DATA1_5 ), .IN2(n14352), .IN3(\U160/DATA1_5 ), 
        .IN4(n14341), .IN5(n9667), .Q(n9664) );
  AO22X1 U1851 ( .IN1(\U150/DATA1_5 ), .IN2(n14331), .IN3(\U155/DATA1_5 ), 
        .IN4(n14314), .Q(n9667) );
  AO221X1 U1852 ( .IN1(n5370), .IN2(n14249), .IN3(\U125/DATA1_4 ), .IN4(n14194), .IN5(n9668), .Q(n13192) );
  AO222X1 U1853 ( .IN1(\U130/DATA1_4 ), .IN2(n14409), .IN3(n14399), .IN4(n9669), .IN5(\U135/DATA1_4 ), .IN6(n14388), .Q(n9668) );
  OR2X1 U1854 ( .IN1(n9670), .IN2(n9671), .Q(n9669) );
  AO221X1 U1855 ( .IN1(\U165/DATA1_4 ), .IN2(n14383), .IN3(\U170/DATA1_4 ), 
        .IN4(n14371), .IN5(n9672), .Q(n9671) );
  AO22X1 U1856 ( .IN1(\U140/DATA1_4 ), .IN2(n14256), .IN3(\U170/DATA2_4 ), 
        .IN4(n14358), .Q(n9672) );
  AO221X1 U1857 ( .IN1(\U145/DATA1_4 ), .IN2(n14352), .IN3(\U160/DATA1_4 ), 
        .IN4(n14341), .IN5(n9673), .Q(n9670) );
  AO22X1 U1858 ( .IN1(\U150/DATA1_4 ), .IN2(n14331), .IN3(\U155/DATA1_4 ), 
        .IN4(n14318), .Q(n9673) );
  AO221X1 U1859 ( .IN1(n5369), .IN2(n14249), .IN3(\U125/DATA1_3 ), .IN4(n14194), .IN5(n9674), .Q(n13193) );
  AO222X1 U1860 ( .IN1(\U130/DATA1_3 ), .IN2(n14409), .IN3(n14399), .IN4(n9675), .IN5(\U135/DATA1_3 ), .IN6(n14388), .Q(n9674) );
  OR2X1 U1861 ( .IN1(n9676), .IN2(n9677), .Q(n9675) );
  AO221X1 U1862 ( .IN1(\U165/DATA1_3 ), .IN2(n14383), .IN3(\U170/DATA1_3 ), 
        .IN4(n14371), .IN5(n9678), .Q(n9677) );
  AO22X1 U1863 ( .IN1(\U140/DATA1_3 ), .IN2(n14186), .IN3(\U170/DATA2_3 ), 
        .IN4(n14358), .Q(n9678) );
  AO221X1 U1864 ( .IN1(\U145/DATA1_3 ), .IN2(n14352), .IN3(\U160/DATA1_3 ), 
        .IN4(n14341), .IN5(n9679), .Q(n9676) );
  AO22X1 U1865 ( .IN1(\U150/DATA1_3 ), .IN2(n14331), .IN3(\U155/DATA1_3 ), 
        .IN4(n14313), .Q(n9679) );
  AO221X1 U1866 ( .IN1(n5368), .IN2(n14249), .IN3(\U125/DATA1_2 ), .IN4(n14194), .IN5(n9680), .Q(n13194) );
  AO222X1 U1867 ( .IN1(\U130/DATA1_2 ), .IN2(n14409), .IN3(n14399), .IN4(n9681), .IN5(\U135/DATA1_2 ), .IN6(n14388), .Q(n9680) );
  OR2X1 U1868 ( .IN1(n9682), .IN2(n9683), .Q(n9681) );
  AO221X1 U1869 ( .IN1(\U165/DATA1_2 ), .IN2(n14383), .IN3(\U170/DATA1_2 ), 
        .IN4(n14371), .IN5(n9684), .Q(n9683) );
  AO22X1 U1870 ( .IN1(\U140/DATA1_2 ), .IN2(n14257), .IN3(\U170/DATA2_2 ), 
        .IN4(n14358), .Q(n9684) );
  AO221X1 U1871 ( .IN1(\U145/DATA1_2 ), .IN2(n14352), .IN3(\U160/DATA1_2 ), 
        .IN4(n14341), .IN5(n9685), .Q(n9682) );
  AO22X1 U1872 ( .IN1(\U150/DATA1_2 ), .IN2(n14331), .IN3(\U155/DATA1_2 ), 
        .IN4(n14317), .Q(n9685) );
  AO221X1 U1873 ( .IN1(n5367), .IN2(n14249), .IN3(\U125/DATA1_1 ), .IN4(n14194), .IN5(n9686), .Q(n13195) );
  AO222X1 U1874 ( .IN1(\U130/DATA1_1 ), .IN2(n14409), .IN3(n14399), .IN4(n9687), .IN5(\U135/DATA1_1 ), .IN6(n14388), .Q(n9686) );
  OR2X1 U1875 ( .IN1(n9688), .IN2(n9689), .Q(n9687) );
  AO221X1 U1876 ( .IN1(p___constant_11x11xf32_8_2[1]), .IN2(n14383), .IN3(
        p___constant_11x11xf32_8_1[1]), .IN4(n14371), .IN5(n9690), .Q(n9689)
         );
  AO22X1 U1877 ( .IN1(\U140/DATA1_1 ), .IN2(n14192), .IN3(
        p___constant_11x11xf32_8_0[1]), .IN4(n14358), .Q(n9690) );
  AO221X1 U1878 ( .IN1(p___constant_11x11xf32_8_6[1]), .IN2(n14352), .IN3(
        p___constant_11x11xf32_8_3[1]), .IN4(n14341), .IN5(n9691), .Q(n9688)
         );
  AO22X1 U1879 ( .IN1(p___constant_11x11xf32_8_5[1]), .IN2(n14331), .IN3(
        p___constant_11x11xf32_8_4[1]), .IN4(n14317), .Q(n9691) );
  AO221X1 U1880 ( .IN1(n5366), .IN2(n14237), .IN3(\U125/DATA1_0 ), .IN4(n14194), .IN5(n9692), .Q(n13196) );
  AO222X1 U1881 ( .IN1(\U130/DATA1_0 ), .IN2(n14409), .IN3(n14399), .IN4(n9693), .IN5(\U135/DATA1_0 ), .IN6(n14388), .Q(n9692) );
  OR2X1 U1882 ( .IN1(n9694), .IN2(n9695), .Q(n9693) );
  AO221X1 U1883 ( .IN1(p___constant_11x11xf32_8_2[0]), .IN2(n14383), .IN3(
        p___constant_11x11xf32_8_1[0]), .IN4(n14371), .IN5(n9696), .Q(n9695)
         );
  AO22X1 U1884 ( .IN1(\U140/DATA1_0 ), .IN2(n14186), .IN3(
        p___constant_11x11xf32_8_0[0]), .IN4(n14358), .Q(n9696) );
  AO221X1 U1885 ( .IN1(p___constant_11x11xf32_8_6[0]), .IN2(n14352), .IN3(
        p___constant_11x11xf32_8_3[0]), .IN4(n14341), .IN5(n9697), .Q(n9694)
         );
  AO22X1 U1886 ( .IN1(p___constant_11x11xf32_8_5[0]), .IN2(n14331), .IN3(
        p___constant_11x11xf32_8_4[0]), .IN4(n14319), .Q(n9697) );
  AO21X1 U1887 ( .IN1(n14240), .IN2(n13763), .IN3(n9529), .Q(n13197) );
  AO21X1 U1888 ( .IN1(n14240), .IN2(n13895), .IN3(n9531), .Q(n13198) );
  AO21X1 U1889 ( .IN1(n14240), .IN2(n14075), .IN3(n9533), .Q(n13199) );
  AO21X1 U1891 ( .IN1(n5386), .IN2(n14243), .IN3(n9534), .Q(n13200) );
  AO21X1 U1892 ( .IN1(n5385), .IN2(n14243), .IN3(n9535), .Q(n13201) );
  AO21X1 U1893 ( .IN1(n5384), .IN2(n14244), .IN3(n9536), .Q(n13202) );
  AO21X1 U1894 ( .IN1(n5383), .IN2(n14243), .IN3(n9537), .Q(n13203) );
  AO21X1 U1895 ( .IN1(n5382), .IN2(n14243), .IN3(n9538), .Q(n13204) );
  AO21X1 U1896 ( .IN1(n5381), .IN2(n14243), .IN3(n9540), .Q(n13205) );
  AO21X1 U1897 ( .IN1(n5380), .IN2(n14243), .IN3(n9542), .Q(n13206) );
  AO21X1 U1898 ( .IN1(n5379), .IN2(n14243), .IN3(n9544), .Q(n13207) );
  AO221X1 U1900 ( .IN1(n14238), .IN2(n13915), .IN3(\U178/DATA1_11 ), .IN4(
        n14194), .IN5(n9702), .Q(n13209) );
  AO222X1 U1901 ( .IN1(\U183/DATA1_11 ), .IN2(n14409), .IN3(n14400), .IN4(
        n9703), .IN5(\U188/DATA1_11 ), .IN6(n14389), .Q(n9702) );
  OR2X1 U1902 ( .IN1(n9704), .IN2(n9705), .Q(n9703) );
  AO221X1 U1903 ( .IN1(\U218/DATA1_11 ), .IN2(n14382), .IN3(\U223/DATA1_11 ), 
        .IN4(n14370), .IN5(n9706), .Q(n9705) );
  AO22X1 U1904 ( .IN1(\U193/DATA1_11 ), .IN2(n14914), .IN3(\U223/DATA2_11 ), 
        .IN4(n14358), .Q(n9706) );
  AO221X1 U1905 ( .IN1(\U198/DATA1_11 ), .IN2(n14351), .IN3(\U213/DATA1_11 ), 
        .IN4(n14340), .IN5(n9707), .Q(n9704) );
  AO22X1 U1906 ( .IN1(\U203/DATA1_11 ), .IN2(n14330), .IN3(\U208/DATA1_11 ), 
        .IN4(n14320), .Q(n9707) );
  AO221X1 U1908 ( .IN1(n14236), .IN2(n13905), .IN3(\U178/DATA1_10 ), .IN4(
        n14194), .IN5(n9709), .Q(n13210) );
  AO222X1 U1909 ( .IN1(\U183/DATA1_10 ), .IN2(n14409), .IN3(n14400), .IN4(
        n9710), .IN5(\U188/DATA1_10 ), .IN6(n14389), .Q(n9709) );
  OR2X1 U1910 ( .IN1(n9711), .IN2(n9712), .Q(n9710) );
  AO221X1 U1911 ( .IN1(\U218/DATA1_10 ), .IN2(n14382), .IN3(\U223/DATA1_10 ), 
        .IN4(n14370), .IN5(n9713), .Q(n9712) );
  AO22X1 U1912 ( .IN1(\U193/DATA1_10 ), .IN2(n14191), .IN3(\U223/DATA2_10 ), 
        .IN4(n14358), .Q(n9713) );
  AO221X1 U1913 ( .IN1(\U198/DATA1_10 ), .IN2(n14351), .IN3(\U213/DATA1_10 ), 
        .IN4(n14340), .IN5(n9714), .Q(n9711) );
  AO22X1 U1914 ( .IN1(\U203/DATA1_10 ), .IN2(n14330), .IN3(\U208/DATA1_10 ), 
        .IN4(n14320), .Q(n9714) );
  AO221X1 U1915 ( .IN1(n14238), .IN2(n14047), .IN3(\U178/DATA1_9 ), .IN4(
        n14194), .IN5(n9716), .Q(n13211) );
  AO222X1 U1916 ( .IN1(\U183/DATA1_9 ), .IN2(n14409), .IN3(n14400), .IN4(n9717), .IN5(\U188/DATA1_9 ), .IN6(n14389), .Q(n9716) );
  OR2X1 U1917 ( .IN1(n9718), .IN2(n9719), .Q(n9717) );
  AO221X1 U1918 ( .IN1(\U218/DATA1_9 ), .IN2(n14382), .IN3(\U223/DATA1_9 ), 
        .IN4(n14370), .IN5(n9720), .Q(n9719) );
  AO22X1 U1919 ( .IN1(\U193/DATA1_9 ), .IN2(n14254), .IN3(\U223/DATA2_9 ), 
        .IN4(n14358), .Q(n9720) );
  AO221X1 U1920 ( .IN1(\U198/DATA1_9 ), .IN2(n14351), .IN3(\U213/DATA1_9 ), 
        .IN4(n14340), .IN5(n9721), .Q(n9718) );
  AO22X1 U1921 ( .IN1(\U203/DATA1_9 ), .IN2(n14330), .IN3(\U208/DATA1_9 ), 
        .IN4(n14320), .Q(n9721) );
  AO221X1 U1923 ( .IN1(n5446), .IN2(n14905), .IN3(\U178/DATA1_8 ), .IN4(n14194), .IN5(n9722), .Q(n13212) );
  AO222X1 U1924 ( .IN1(\U183/DATA1_8 ), .IN2(n14409), .IN3(n14400), .IN4(n9723), .IN5(\U188/DATA1_8 ), .IN6(n14389), .Q(n9722) );
  OR2X1 U1925 ( .IN1(n9724), .IN2(n9725), .Q(n9723) );
  AO221X1 U1926 ( .IN1(\U218/DATA1_8 ), .IN2(n14382), .IN3(\U223/DATA1_8 ), 
        .IN4(n14370), .IN5(n9726), .Q(n9725) );
  AO22X1 U1927 ( .IN1(\U193/DATA1_8 ), .IN2(n14257), .IN3(\U223/DATA2_8 ), 
        .IN4(n14358), .Q(n9726) );
  AO221X1 U1928 ( .IN1(\U198/DATA1_8 ), .IN2(n14351), .IN3(\U213/DATA1_8 ), 
        .IN4(n14340), .IN5(n9727), .Q(n9724) );
  AO22X1 U1929 ( .IN1(\U203/DATA1_8 ), .IN2(n14330), .IN3(\U208/DATA1_8 ), 
        .IN4(n14320), .Q(n9727) );
  AO221X1 U1930 ( .IN1(n5445), .IN2(n14246), .IN3(\U178/DATA1_7 ), .IN4(n14194), .IN5(n9728), .Q(n13213) );
  AO222X1 U1931 ( .IN1(\U183/DATA1_7 ), .IN2(n14409), .IN3(n14400), .IN4(n9729), .IN5(\U188/DATA1_7 ), .IN6(n14389), .Q(n9728) );
  OR2X1 U1932 ( .IN1(n9730), .IN2(n9731), .Q(n9729) );
  AO221X1 U1933 ( .IN1(\U218/DATA1_7 ), .IN2(n14382), .IN3(\U223/DATA1_7 ), 
        .IN4(n14370), .IN5(n9732), .Q(n9731) );
  AO22X1 U1934 ( .IN1(\U193/DATA1_7 ), .IN2(n14914), .IN3(\U223/DATA2_7 ), 
        .IN4(n14361), .Q(n9732) );
  AO221X1 U1935 ( .IN1(\U198/DATA1_7 ), .IN2(n14351), .IN3(\U213/DATA1_7 ), 
        .IN4(n14340), .IN5(n9733), .Q(n9730) );
  AO22X1 U1936 ( .IN1(\U203/DATA1_7 ), .IN2(n14330), .IN3(\U208/DATA1_7 ), 
        .IN4(n14320), .Q(n9733) );
  AO221X1 U1937 ( .IN1(n5444), .IN2(n14250), .IN3(
        p___constant_11x11xf32_7_10[6]), .IN4(n14195), .IN5(n9734), .Q(n13214)
         );
  AO222X1 U1938 ( .IN1(p___constant_11x11xf32_7_9[6]), .IN2(n14409), .IN3(
        n14400), .IN4(n9735), .IN5(p___constant_11x11xf32_7_8[6]), .IN6(n14389), .Q(n9734) );
  OR2X1 U1939 ( .IN1(n9736), .IN2(n9737), .Q(n9735) );
  AO221X1 U1940 ( .IN1(\U218/DATA1_6 ), .IN2(n14382), .IN3(\U223/DATA1_6 ), 
        .IN4(n14370), .IN5(n9738), .Q(n9737) );
  AO22X1 U1941 ( .IN1(p___constant_11x11xf32_7_7[6]), .IN2(n14914), .IN3(
        \U223/DATA2_6 ), .IN4(n14360), .Q(n9738) );
  AO221X1 U1942 ( .IN1(p___constant_11x11xf32_7_6[6]), .IN2(n14351), .IN3(
        \U213/DATA1_6 ), .IN4(n14340), .IN5(n9739), .Q(n9736) );
  AO22X1 U1943 ( .IN1(p___constant_11x11xf32_7_5[6]), .IN2(n14330), .IN3(
        \U208/DATA1_6 ), .IN4(n14320), .Q(n9739) );
  AO221X1 U1944 ( .IN1(n5443), .IN2(n14234), .IN3(
        p___constant_11x11xf32_7_10[5]), .IN4(n14195), .IN5(n9740), .Q(n13215)
         );
  AO222X1 U1945 ( .IN1(p___constant_11x11xf32_7_9[5]), .IN2(n14409), .IN3(
        n14400), .IN4(n9741), .IN5(p___constant_11x11xf32_7_8[5]), .IN6(n14389), .Q(n9740) );
  OR2X1 U1946 ( .IN1(n9742), .IN2(n9743), .Q(n9741) );
  AO221X1 U1947 ( .IN1(p___constant_11x11xf32_7_2[5]), .IN2(n14382), .IN3(
        p___constant_11x11xf32_7_1[5]), .IN4(n14370), .IN5(n9744), .Q(n9743)
         );
  AO22X1 U1948 ( .IN1(p___constant_11x11xf32_7_7[5]), .IN2(n14191), .IN3(
        p___constant_11x11xf32_7_0[5]), .IN4(n14362), .Q(n9744) );
  AO221X1 U1949 ( .IN1(p___constant_11x11xf32_7_6[5]), .IN2(n14351), .IN3(
        p___constant_11x11xf32_7_3[5]), .IN4(n14340), .IN5(n9745), .Q(n9742)
         );
  AO22X1 U1950 ( .IN1(p___constant_11x11xf32_7_5[5]), .IN2(n14330), .IN3(
        p___constant_11x11xf32_7_4[5]), .IN4(n14320), .Q(n9745) );
  AO221X1 U1951 ( .IN1(n5442), .IN2(n14242), .IN3(
        p___constant_11x11xf32_7_10[4]), .IN4(n14195), .IN5(n9746), .Q(n13216)
         );
  AO222X1 U1952 ( .IN1(p___constant_11x11xf32_7_9[4]), .IN2(n14409), .IN3(
        n14400), .IN4(n9747), .IN5(p___constant_11x11xf32_7_8[4]), .IN6(n14389), .Q(n9746) );
  OR2X1 U1953 ( .IN1(n9748), .IN2(n9749), .Q(n9747) );
  AO221X1 U1954 ( .IN1(p___constant_11x11xf32_7_2[4]), .IN2(n14382), .IN3(
        p___constant_11x11xf32_7_1[4]), .IN4(n14370), .IN5(n9750), .Q(n9749)
         );
  AO22X1 U1955 ( .IN1(p___constant_11x11xf32_7_7[4]), .IN2(n14914), .IN3(
        p___constant_11x11xf32_7_0[4]), .IN4(n14362), .Q(n9750) );
  AO221X1 U1956 ( .IN1(p___constant_11x11xf32_7_6[4]), .IN2(n14351), .IN3(
        p___constant_11x11xf32_7_3[4]), .IN4(n14340), .IN5(n9751), .Q(n9748)
         );
  AO22X1 U1957 ( .IN1(p___constant_11x11xf32_7_5[4]), .IN2(n14330), .IN3(
        p___constant_11x11xf32_7_4[4]), .IN4(n14320), .Q(n9751) );
  AO221X1 U1958 ( .IN1(n5441), .IN2(n14247), .IN3(
        p___constant_11x11xf32_7_10[3]), .IN4(n14195), .IN5(n9752), .Q(n13217)
         );
  AO222X1 U1959 ( .IN1(p___constant_11x11xf32_7_9[3]), .IN2(n14409), .IN3(
        n14400), .IN4(n9753), .IN5(p___constant_11x11xf32_7_8[3]), .IN6(n14389), .Q(n9752) );
  OR2X1 U1960 ( .IN1(n9754), .IN2(n9755), .Q(n9753) );
  AO221X1 U1961 ( .IN1(p___constant_11x11xf32_7_2[3]), .IN2(n14382), .IN3(
        p___constant_11x11xf32_7_1[3]), .IN4(n14370), .IN5(n9756), .Q(n9755)
         );
  AO22X1 U1962 ( .IN1(p___constant_11x11xf32_7_7[3]), .IN2(n14186), .IN3(
        p___constant_11x11xf32_7_0[3]), .IN4(n14362), .Q(n9756) );
  AO221X1 U1963 ( .IN1(p___constant_11x11xf32_7_6[3]), .IN2(n14351), .IN3(
        p___constant_11x11xf32_7_3[3]), .IN4(n14340), .IN5(n9757), .Q(n9754)
         );
  AO22X1 U1964 ( .IN1(p___constant_11x11xf32_7_5[3]), .IN2(n14330), .IN3(
        p___constant_11x11xf32_7_4[3]), .IN4(n14320), .Q(n9757) );
  AO221X1 U1965 ( .IN1(n5440), .IN2(n14246), .IN3(
        p___constant_11x11xf32_7_10[2]), .IN4(n14195), .IN5(n9758), .Q(n13218)
         );
  AO222X1 U1966 ( .IN1(p___constant_11x11xf32_7_9[2]), .IN2(n14409), .IN3(
        n14400), .IN4(n9759), .IN5(p___constant_11x11xf32_7_8[2]), .IN6(n14389), .Q(n9758) );
  OR2X1 U1967 ( .IN1(n9760), .IN2(n9761), .Q(n9759) );
  AO221X1 U1968 ( .IN1(p___constant_11x11xf32_7_2[2]), .IN2(n14382), .IN3(
        p___constant_11x11xf32_7_1[2]), .IN4(n14370), .IN5(n9762), .Q(n9761)
         );
  AO22X1 U1969 ( .IN1(p___constant_11x11xf32_7_7[2]), .IN2(n14186), .IN3(
        p___constant_11x11xf32_7_0[2]), .IN4(n14356), .Q(n9762) );
  AO221X1 U1970 ( .IN1(p___constant_11x11xf32_7_6[2]), .IN2(n14351), .IN3(
        p___constant_11x11xf32_7_3[2]), .IN4(n14340), .IN5(n9763), .Q(n9760)
         );
  AO22X1 U1971 ( .IN1(p___constant_11x11xf32_7_5[2]), .IN2(n14330), .IN3(
        p___constant_11x11xf32_7_4[2]), .IN4(n14320), .Q(n9763) );
  AO221X1 U1972 ( .IN1(n5439), .IN2(n14243), .IN3(
        p___constant_11x11xf32_7_10[1]), .IN4(n14195), .IN5(n9764), .Q(n13219)
         );
  AO222X1 U1973 ( .IN1(p___constant_11x11xf32_7_9[1]), .IN2(n14406), .IN3(
        n14400), .IN4(n9765), .IN5(p___constant_11x11xf32_7_8[1]), .IN6(n14389), .Q(n9764) );
  OR2X1 U1974 ( .IN1(n9766), .IN2(n9767), .Q(n9765) );
  AO221X1 U1975 ( .IN1(p___constant_11x11xf32_7_2[1]), .IN2(n14382), .IN3(
        p___constant_11x11xf32_7_1[1]), .IN4(n14370), .IN5(n9768), .Q(n9767)
         );
  AO22X1 U1976 ( .IN1(p___constant_11x11xf32_7_7[1]), .IN2(n14254), .IN3(
        p___constant_11x11xf32_7_0[1]), .IN4(n14360), .Q(n9768) );
  AO221X1 U1977 ( .IN1(p___constant_11x11xf32_7_6[1]), .IN2(n14351), .IN3(
        p___constant_11x11xf32_7_3[1]), .IN4(n14340), .IN5(n9769), .Q(n9766)
         );
  AO22X1 U1978 ( .IN1(p___constant_11x11xf32_7_5[1]), .IN2(n14330), .IN3(
        p___constant_11x11xf32_7_4[1]), .IN4(n14320), .Q(n9769) );
  AO221X1 U1979 ( .IN1(n5438), .IN2(n14241), .IN3(
        p___constant_11x11xf32_7_10[0]), .IN4(n14195), .IN5(n9770), .Q(n13220)
         );
  AO222X1 U1980 ( .IN1(p___constant_11x11xf32_7_9[0]), .IN2(n14407), .IN3(
        n14400), .IN4(n9771), .IN5(p___constant_11x11xf32_7_8[0]), .IN6(n14389), .Q(n9770) );
  OR2X1 U1981 ( .IN1(n9772), .IN2(n9773), .Q(n9771) );
  AO221X1 U1982 ( .IN1(p___constant_11x11xf32_7_2[0]), .IN2(n14382), .IN3(
        p___constant_11x11xf32_7_1[0]), .IN4(n14370), .IN5(n9774), .Q(n9773)
         );
  AO22X1 U1983 ( .IN1(p___constant_11x11xf32_7_7[0]), .IN2(n14914), .IN3(
        p___constant_11x11xf32_7_0[0]), .IN4(n14363), .Q(n9774) );
  AO221X1 U1984 ( .IN1(p___constant_11x11xf32_7_6[0]), .IN2(n14351), .IN3(
        p___constant_11x11xf32_7_3[0]), .IN4(n14340), .IN5(n9775), .Q(n9772)
         );
  AO22X1 U1985 ( .IN1(p___constant_11x11xf32_7_5[0]), .IN2(n14330), .IN3(
        p___constant_11x11xf32_7_4[0]), .IN4(n14320), .Q(n9775) );
  AO21X1 U1986 ( .IN1(n14240), .IN2(n13762), .IN3(n9529), .Q(n13221) );
  AO21X1 U1987 ( .IN1(n14240), .IN2(n13615), .IN3(n9531), .Q(n13222) );
  AO21X1 U1988 ( .IN1(n14241), .IN2(n14074), .IN3(n9533), .Q(n13223) );
  AO21X1 U1990 ( .IN1(n5458), .IN2(n14243), .IN3(n9534), .Q(n13224) );
  AO21X1 U1991 ( .IN1(n5457), .IN2(n14243), .IN3(n9535), .Q(n13225) );
  AO21X1 U1992 ( .IN1(n5456), .IN2(n14243), .IN3(n9536), .Q(n13226) );
  AO21X1 U1993 ( .IN1(n5455), .IN2(n14243), .IN3(n9537), .Q(n13227) );
  AO21X1 U1994 ( .IN1(n5454), .IN2(n14242), .IN3(n9538), .Q(n13228) );
  AO21X1 U1995 ( .IN1(n5453), .IN2(n14242), .IN3(n9540), .Q(n13229) );
  AO21X1 U1996 ( .IN1(n5452), .IN2(n14242), .IN3(n9542), .Q(n13230) );
  AO21X1 U1997 ( .IN1(n5451), .IN2(n14242), .IN3(n9544), .Q(n13231) );
  AO221X1 U1999 ( .IN1(n14238), .IN2(n13914), .IN3(\U234/DATA1_11 ), .IN4(
        n14195), .IN5(n9780), .Q(n13233) );
  AO222X1 U2000 ( .IN1(\U239/DATA1_11 ), .IN2(n14408), .IN3(n14401), .IN4(
        n9781), .IN5(\U244/DATA1_11 ), .IN6(n14391), .Q(n9780) );
  OR2X1 U2001 ( .IN1(n9782), .IN2(n9783), .Q(n9781) );
  AO221X1 U2002 ( .IN1(\U274/DATA1_11 ), .IN2(n14381), .IN3(\U279/DATA1_11 ), 
        .IN4(n14369), .IN5(n9784), .Q(n9783) );
  AO22X1 U2003 ( .IN1(\U249/DATA1_11 ), .IN2(n14189), .IN3(\U279/DATA2_11 ), 
        .IN4(n14362), .Q(n9784) );
  AO221X1 U2004 ( .IN1(\U254/DATA1_11 ), .IN2(n14350), .IN3(\U269/DATA1_11 ), 
        .IN4(n14339), .IN5(n9785), .Q(n9782) );
  AO22X1 U2005 ( .IN1(p___constant_11x11xf32_6_5[11]), .IN2(n14329), .IN3(
        \U264/DATA1_11 ), .IN4(n14319), .Q(n9785) );
  AO221X1 U2007 ( .IN1(n14237), .IN2(n13904), .IN3(\U234/DATA1_10 ), .IN4(
        n14195), .IN5(n9787), .Q(n13234) );
  AO222X1 U2008 ( .IN1(\U239/DATA1_10 ), .IN2(n14410), .IN3(n14401), .IN4(
        n9788), .IN5(\U244/DATA1_10 ), .IN6(n14386), .Q(n9787) );
  OR2X1 U2009 ( .IN1(n9789), .IN2(n9790), .Q(n9788) );
  AO221X1 U2010 ( .IN1(\U274/DATA1_10 ), .IN2(n14381), .IN3(\U279/DATA1_10 ), 
        .IN4(n14369), .IN5(n9791), .Q(n9790) );
  AO22X1 U2011 ( .IN1(\U249/DATA1_10 ), .IN2(n14191), .IN3(\U279/DATA2_10 ), 
        .IN4(n14363), .Q(n9791) );
  AO221X1 U2012 ( .IN1(\U254/DATA1_10 ), .IN2(n14350), .IN3(\U269/DATA1_10 ), 
        .IN4(n14339), .IN5(n9792), .Q(n9789) );
  AO22X1 U2013 ( .IN1(p___constant_11x11xf32_6_5[10]), .IN2(n14329), .IN3(
        \U264/DATA1_10 ), .IN4(n14319), .Q(n9792) );
  AO221X1 U2014 ( .IN1(n14238), .IN2(n14046), .IN3(\U234/DATA1_9 ), .IN4(
        n14195), .IN5(n9794), .Q(n13235) );
  AO222X1 U2015 ( .IN1(\U239/DATA1_9 ), .IN2(n14409), .IN3(n14401), .IN4(n9795), .IN5(\U244/DATA1_9 ), .IN6(n14387), .Q(n9794) );
  OR2X1 U2016 ( .IN1(n9796), .IN2(n9797), .Q(n9795) );
  AO221X1 U2017 ( .IN1(\U274/DATA1_9 ), .IN2(n14381), .IN3(\U279/DATA1_9 ), 
        .IN4(n14369), .IN5(n9798), .Q(n9797) );
  AO22X1 U2018 ( .IN1(\U249/DATA1_9 ), .IN2(n14190), .IN3(\U279/DATA2_9 ), 
        .IN4(n14361), .Q(n9798) );
  AO221X1 U2019 ( .IN1(\U254/DATA1_9 ), .IN2(n14350), .IN3(\U269/DATA1_9 ), 
        .IN4(n14339), .IN5(n9799), .Q(n9796) );
  AO22X1 U2020 ( .IN1(p___constant_11x11xf32_6_5[9]), .IN2(n14329), .IN3(
        \U264/DATA1_9 ), .IN4(n14319), .Q(n9799) );
  AO221X1 U2022 ( .IN1(n5518), .IN2(n14236), .IN3(\U234/DATA1_8 ), .IN4(n14195), .IN5(n9800), .Q(n13236) );
  AO222X1 U2023 ( .IN1(\U239/DATA1_8 ), .IN2(n14406), .IN3(n14401), .IN4(n9801), .IN5(\U244/DATA1_8 ), .IN6(n14388), .Q(n9800) );
  OR2X1 U2024 ( .IN1(n9802), .IN2(n9803), .Q(n9801) );
  AO221X1 U2025 ( .IN1(\U274/DATA1_8 ), .IN2(n14381), .IN3(\U279/DATA1_8 ), 
        .IN4(n14369), .IN5(n9804), .Q(n9803) );
  AO22X1 U2026 ( .IN1(\U249/DATA1_8 ), .IN2(n14193), .IN3(\U279/DATA2_8 ), 
        .IN4(n14357), .Q(n9804) );
  AO221X1 U2027 ( .IN1(\U254/DATA1_8 ), .IN2(n14350), .IN3(\U269/DATA1_8 ), 
        .IN4(n14339), .IN5(n9805), .Q(n9802) );
  AO22X1 U2028 ( .IN1(p___constant_11x11xf32_6_5[8]), .IN2(n14329), .IN3(
        \U264/DATA1_8 ), .IN4(n14319), .Q(n9805) );
  AO221X1 U2029 ( .IN1(n5517), .IN2(n14240), .IN3(\U234/DATA1_7 ), .IN4(n14195), .IN5(n9806), .Q(n13237) );
  AO222X1 U2030 ( .IN1(\U239/DATA1_7 ), .IN2(n14413), .IN3(n14401), .IN4(n9807), .IN5(\U244/DATA1_7 ), .IN6(n14393), .Q(n9806) );
  OR2X1 U2031 ( .IN1(n9808), .IN2(n9809), .Q(n9807) );
  AO221X1 U2032 ( .IN1(\U274/DATA1_7 ), .IN2(n14381), .IN3(\U279/DATA1_7 ), 
        .IN4(n14369), .IN5(n9810), .Q(n9809) );
  AO22X1 U2033 ( .IN1(\U249/DATA1_7 ), .IN2(n14255), .IN3(\U279/DATA2_7 ), 
        .IN4(n14360), .Q(n9810) );
  AO221X1 U2034 ( .IN1(\U254/DATA1_7 ), .IN2(n14350), .IN3(\U269/DATA1_7 ), 
        .IN4(n14339), .IN5(n9811), .Q(n9808) );
  AO22X1 U2035 ( .IN1(p___constant_11x11xf32_6_5[7]), .IN2(n14329), .IN3(
        \U264/DATA1_7 ), .IN4(n14319), .Q(n9811) );
  AO221X1 U2036 ( .IN1(n5516), .IN2(n14235), .IN3(\U234/DATA1_6 ), .IN4(n13736), .IN5(n9812), .Q(n13238) );
  AO222X1 U2037 ( .IN1(\U239/DATA1_6 ), .IN2(n14406), .IN3(n14401), .IN4(n9813), .IN5(\U244/DATA1_6 ), .IN6(n14387), .Q(n9812) );
  OR2X1 U2038 ( .IN1(n9814), .IN2(n9815), .Q(n9813) );
  AO221X1 U2039 ( .IN1(\U274/DATA1_6 ), .IN2(n14381), .IN3(\U279/DATA1_6 ), 
        .IN4(n14369), .IN5(n9816), .Q(n9815) );
  AO22X1 U2040 ( .IN1(\U249/DATA1_6 ), .IN2(n14255), .IN3(\U279/DATA2_6 ), 
        .IN4(n14360), .Q(n9816) );
  AO221X1 U2041 ( .IN1(\U254/DATA1_6 ), .IN2(n14350), .IN3(\U269/DATA1_6 ), 
        .IN4(n14339), .IN5(n9817), .Q(n9814) );
  AO22X1 U2042 ( .IN1(p___constant_11x11xf32_6_5[6]), .IN2(n14329), .IN3(
        \U264/DATA1_6 ), .IN4(n14319), .Q(n9817) );
  AO221X1 U2043 ( .IN1(n5515), .IN2(n14241), .IN3(\U234/DATA1_5 ), .IN4(n13736), .IN5(n9818), .Q(n13239) );
  AO222X1 U2044 ( .IN1(\U239/DATA1_5 ), .IN2(n14406), .IN3(n14401), .IN4(n9819), .IN5(\U244/DATA1_5 ), .IN6(n14389), .Q(n9818) );
  OR2X1 U2045 ( .IN1(n9820), .IN2(n9821), .Q(n9819) );
  AO221X1 U2046 ( .IN1(\U274/DATA1_5 ), .IN2(n14381), .IN3(\U279/DATA1_5 ), 
        .IN4(n14369), .IN5(n9822), .Q(n9821) );
  AO22X1 U2047 ( .IN1(\U249/DATA1_5 ), .IN2(n14256), .IN3(\U279/DATA2_5 ), 
        .IN4(n14360), .Q(n9822) );
  AO221X1 U2048 ( .IN1(\U254/DATA1_5 ), .IN2(n14350), .IN3(\U269/DATA1_5 ), 
        .IN4(n14339), .IN5(n9823), .Q(n9820) );
  AO22X1 U2049 ( .IN1(p___constant_11x11xf32_6_5[5]), .IN2(n14329), .IN3(
        \U264/DATA1_5 ), .IN4(n14319), .Q(n9823) );
  AO221X1 U2050 ( .IN1(n5514), .IN2(n14234), .IN3(\U234/DATA1_4 ), .IN4(n13736), .IN5(n9824), .Q(n13240) );
  AO222X1 U2051 ( .IN1(\U239/DATA1_4 ), .IN2(n14406), .IN3(n14401), .IN4(n9825), .IN5(\U244/DATA1_4 ), .IN6(n14391), .Q(n9824) );
  OR2X1 U2052 ( .IN1(n9826), .IN2(n9827), .Q(n9825) );
  AO221X1 U2053 ( .IN1(\U274/DATA1_4 ), .IN2(n14381), .IN3(\U279/DATA1_4 ), 
        .IN4(n14369), .IN5(n9828), .Q(n9827) );
  AO22X1 U2054 ( .IN1(\U249/DATA1_4 ), .IN2(n14255), .IN3(\U279/DATA2_4 ), 
        .IN4(n14359), .Q(n9828) );
  AO221X1 U2055 ( .IN1(\U254/DATA1_4 ), .IN2(n14350), .IN3(\U269/DATA1_4 ), 
        .IN4(n14339), .IN5(n9829), .Q(n9826) );
  AO22X1 U2056 ( .IN1(p___constant_11x11xf32_6_5[4]), .IN2(n14329), .IN3(
        \U264/DATA1_4 ), .IN4(n14319), .Q(n9829) );
  AO221X1 U2057 ( .IN1(n5513), .IN2(n14905), .IN3(\U234/DATA1_3 ), .IN4(n13736), .IN5(n9830), .Q(n13241) );
  AO222X1 U2058 ( .IN1(\U239/DATA1_3 ), .IN2(n14407), .IN3(n14401), .IN4(n9831), .IN5(\U244/DATA1_3 ), .IN6(n14390), .Q(n9830) );
  OR2X1 U2059 ( .IN1(n9832), .IN2(n9833), .Q(n9831) );
  AO221X1 U2060 ( .IN1(\U274/DATA1_3 ), .IN2(n14381), .IN3(\U279/DATA1_3 ), 
        .IN4(n14369), .IN5(n9834), .Q(n9833) );
  AO22X1 U2061 ( .IN1(\U249/DATA1_3 ), .IN2(n14914), .IN3(\U279/DATA2_3 ), 
        .IN4(n14361), .Q(n9834) );
  AO221X1 U2062 ( .IN1(\U254/DATA1_3 ), .IN2(n14350), .IN3(\U269/DATA1_3 ), 
        .IN4(n14339), .IN5(n9835), .Q(n9832) );
  AO22X1 U2063 ( .IN1(p___constant_11x11xf32_6_5[3]), .IN2(n14329), .IN3(
        \U264/DATA1_3 ), .IN4(n14319), .Q(n9835) );
  AO221X1 U2064 ( .IN1(n5512), .IN2(n14905), .IN3(\U234/DATA1_2 ), .IN4(n13736), .IN5(n9836), .Q(n13242) );
  AO222X1 U2065 ( .IN1(\U239/DATA1_2 ), .IN2(n14408), .IN3(n14401), .IN4(n9837), .IN5(p___constant_11x11xf32_6_8[2]), .IN6(n14391), .Q(n9836) );
  OR2X1 U2066 ( .IN1(n9838), .IN2(n9839), .Q(n9837) );
  AO221X1 U2067 ( .IN1(\U274/DATA1_2 ), .IN2(n14381), .IN3(\U279/DATA1_2 ), 
        .IN4(n14369), .IN5(n9840), .Q(n9839) );
  AO22X1 U2068 ( .IN1(\U249/DATA1_2 ), .IN2(n14189), .IN3(\U279/DATA2_2 ), 
        .IN4(n14362), .Q(n9840) );
  AO221X1 U2069 ( .IN1(\U254/DATA1_2 ), .IN2(n14350), .IN3(\U269/DATA1_2 ), 
        .IN4(n14339), .IN5(n9841), .Q(n9838) );
  AO22X1 U2070 ( .IN1(p___constant_11x11xf32_6_5[2]), .IN2(n14329), .IN3(
        \U264/DATA1_2 ), .IN4(n14319), .Q(n9841) );
  AO221X1 U2071 ( .IN1(n5511), .IN2(n14247), .IN3(\U234/DATA1_1 ), .IN4(n13736), .IN5(n9842), .Q(n13243) );
  AO222X1 U2072 ( .IN1(\U239/DATA1_1 ), .IN2(n14406), .IN3(n14401), .IN4(n9843), .IN5(p___constant_11x11xf32_6_8[1]), .IN6(n14392), .Q(n9842) );
  OR2X1 U2073 ( .IN1(n9844), .IN2(n9845), .Q(n9843) );
  AO221X1 U2074 ( .IN1(p___constant_11x11xf32_6_2[1]), .IN2(n14381), .IN3(
        \U279/DATA1_1 ), .IN4(n14369), .IN5(n9846), .Q(n9845) );
  AO22X1 U2075 ( .IN1(p___constant_11x11xf32_6_7[1]), .IN2(n14914), .IN3(
        \U279/DATA2_1 ), .IN4(n14355), .Q(n9846) );
  AO221X1 U2076 ( .IN1(\U254/DATA1_1 ), .IN2(n14350), .IN3(\U269/DATA1_1 ), 
        .IN4(n14339), .IN5(n9847), .Q(n9844) );
  AO22X1 U2077 ( .IN1(p___constant_11x11xf32_6_5[1]), .IN2(n14329), .IN3(
        \U264/DATA1_1 ), .IN4(n14319), .Q(n9847) );
  AO221X1 U2078 ( .IN1(n5510), .IN2(n14241), .IN3(
        p___constant_11x11xf32_6_10[0]), .IN4(n13736), .IN5(n9848), .Q(n13244)
         );
  AO222X1 U2079 ( .IN1(p___constant_11x11xf32_6_9[0]), .IN2(n14408), .IN3(
        n14401), .IN4(n9849), .IN5(p___constant_11x11xf32_6_8[0]), .IN6(n14392), .Q(n9848) );
  OR2X1 U2080 ( .IN1(n9850), .IN2(n9851), .Q(n9849) );
  AO221X1 U2081 ( .IN1(p___constant_11x11xf32_6_2[0]), .IN2(n14381), .IN3(
        p___constant_11x11xf32_6_1[0]), .IN4(n14369), .IN5(n9852), .Q(n9851)
         );
  AO22X1 U2082 ( .IN1(p___constant_11x11xf32_6_7[0]), .IN2(n14254), .IN3(
        p___constant_11x11xf32_6_0[0]), .IN4(n14358), .Q(n9852) );
  AO221X1 U2083 ( .IN1(p___constant_11x11xf32_6_6[0]), .IN2(n14350), .IN3(
        p___constant_11x11xf32_6_3[0]), .IN4(n14339), .IN5(n9853), .Q(n9850)
         );
  AO22X1 U2084 ( .IN1(p___constant_11x11xf32_6_5[0]), .IN2(n14329), .IN3(
        p___constant_11x11xf32_6_4[0]), .IN4(n14319), .Q(n9853) );
  AO21X1 U2085 ( .IN1(n14241), .IN2(n13761), .IN3(n9529), .Q(n13245) );
  AO21X1 U2086 ( .IN1(n14241), .IN2(n13614), .IN3(n9531), .Q(n13246) );
  AO21X1 U2087 ( .IN1(n14241), .IN2(n14073), .IN3(n9533), .Q(n13247) );
  AO21X1 U2089 ( .IN1(n5530), .IN2(n14242), .IN3(n9534), .Q(n13248) );
  AO21X1 U2090 ( .IN1(n5529), .IN2(n14242), .IN3(n9535), .Q(n13249) );
  AO21X1 U2091 ( .IN1(n5528), .IN2(n14242), .IN3(n9536), .Q(n13250) );
  AO21X1 U2092 ( .IN1(n5527), .IN2(n14242), .IN3(n9537), .Q(n13251) );
  AO21X1 U2093 ( .IN1(n5526), .IN2(n14242), .IN3(n9538), .Q(n13252) );
  AO21X1 U2094 ( .IN1(n5525), .IN2(n14241), .IN3(n9540), .Q(n13253) );
  AO21X1 U2095 ( .IN1(n5524), .IN2(n14242), .IN3(n9542), .Q(n13254) );
  AO21X1 U2096 ( .IN1(n5523), .IN2(n14241), .IN3(n9544), .Q(n13255) );
  AO221X1 U2098 ( .IN1(n14237), .IN2(n13913), .IN3(\U287/DATA1_11 ), .IN4(
        n14196), .IN5(n9858), .Q(n13257) );
  AO222X1 U2099 ( .IN1(\U292/DATA1_11 ), .IN2(n14414), .IN3(n14402), .IN4(
        n9859), .IN5(\U297/DATA1_11 ), .IN6(n14392), .Q(n9858) );
  OR2X1 U2100 ( .IN1(n9860), .IN2(n9861), .Q(n9859) );
  AO221X1 U2101 ( .IN1(\U327/DATA1_11 ), .IN2(n14382), .IN3(\U332/DATA1_11 ), 
        .IN4(n14368), .IN5(n9862), .Q(n9861) );
  AO22X1 U2102 ( .IN1(\U302/DATA1_11 ), .IN2(n14193), .IN3(\U332/DATA2_11 ), 
        .IN4(n14355), .Q(n9862) );
  AO221X1 U2103 ( .IN1(\U307/DATA1_11 ), .IN2(n14351), .IN3(\U322/DATA1_11 ), 
        .IN4(n14338), .IN5(n9863), .Q(n9860) );
  AO22X1 U2104 ( .IN1(\U312/DATA1_11 ), .IN2(n14328), .IN3(\U317/DATA1_11 ), 
        .IN4(n14318), .Q(n9863) );
  AO221X1 U2106 ( .IN1(n14237), .IN2(n13903), .IN3(\U287/DATA1_10 ), .IN4(
        n14196), .IN5(n9865), .Q(n13258) );
  AO222X1 U2107 ( .IN1(\U292/DATA1_10 ), .IN2(n14410), .IN3(n14402), .IN4(
        n9866), .IN5(\U297/DATA1_10 ), .IN6(n14393), .Q(n9865) );
  OR2X1 U2108 ( .IN1(n9867), .IN2(n9868), .Q(n9866) );
  AO221X1 U2109 ( .IN1(\U327/DATA1_10 ), .IN2(n14376), .IN3(\U332/DATA1_10 ), 
        .IN4(n14368), .IN5(n9869), .Q(n9868) );
  AO22X1 U2110 ( .IN1(\U302/DATA1_10 ), .IN2(n14186), .IN3(\U332/DATA2_10 ), 
        .IN4(n14356), .Q(n9869) );
  AO221X1 U2111 ( .IN1(\U307/DATA1_10 ), .IN2(n14345), .IN3(\U322/DATA1_10 ), 
        .IN4(n14338), .IN5(n9870), .Q(n9867) );
  AO22X1 U2112 ( .IN1(\U312/DATA1_10 ), .IN2(n14328), .IN3(\U317/DATA1_10 ), 
        .IN4(n14318), .Q(n9870) );
  AO221X1 U2113 ( .IN1(n14236), .IN2(n14045), .IN3(\U287/DATA1_9 ), .IN4(
        n14196), .IN5(n9872), .Q(n13259) );
  AO222X1 U2114 ( .IN1(\U292/DATA1_9 ), .IN2(n14410), .IN3(n14402), .IN4(n9873), .IN5(\U297/DATA1_9 ), .IN6(n14394), .Q(n9872) );
  OR2X1 U2115 ( .IN1(n9874), .IN2(n9875), .Q(n9873) );
  AO221X1 U2116 ( .IN1(\U327/DATA1_9 ), .IN2(n14381), .IN3(\U332/DATA1_9 ), 
        .IN4(n14368), .IN5(n9876), .Q(n9875) );
  AO22X1 U2117 ( .IN1(\U302/DATA1_9 ), .IN2(n14255), .IN3(\U332/DATA2_9 ), 
        .IN4(n14362), .Q(n9876) );
  AO221X1 U2118 ( .IN1(\U307/DATA1_9 ), .IN2(n14350), .IN3(\U322/DATA1_9 ), 
        .IN4(n14338), .IN5(n9877), .Q(n9874) );
  AO22X1 U2119 ( .IN1(\U312/DATA1_9 ), .IN2(n14328), .IN3(\U317/DATA1_9 ), 
        .IN4(n14318), .Q(n9877) );
  AO221X1 U2121 ( .IN1(n5590), .IN2(n14247), .IN3(\U287/DATA1_8 ), .IN4(n14196), .IN5(n9878), .Q(n13260) );
  AO222X1 U2122 ( .IN1(\U292/DATA1_8 ), .IN2(n14410), .IN3(n14402), .IN4(n9879), .IN5(\U297/DATA1_8 ), .IN6(n14386), .Q(n9878) );
  OR2X1 U2123 ( .IN1(n9880), .IN2(n9881), .Q(n9879) );
  AO221X1 U2124 ( .IN1(\U327/DATA1_8 ), .IN2(n14380), .IN3(\U332/DATA1_8 ), 
        .IN4(n14368), .IN5(n9882), .Q(n9881) );
  AO22X1 U2125 ( .IN1(\U302/DATA1_8 ), .IN2(n14189), .IN3(\U332/DATA2_8 ), 
        .IN4(n14363), .Q(n9882) );
  AO221X1 U2126 ( .IN1(\U307/DATA1_8 ), .IN2(n14353), .IN3(\U322/DATA1_8 ), 
        .IN4(n14338), .IN5(n9883), .Q(n9880) );
  AO22X1 U2127 ( .IN1(\U312/DATA1_8 ), .IN2(n14328), .IN3(\U317/DATA1_8 ), 
        .IN4(n14318), .Q(n9883) );
  AO221X1 U2128 ( .IN1(n5589), .IN2(n14247), .IN3(\U287/DATA1_7 ), .IN4(n14196), .IN5(n9884), .Q(n13261) );
  AO222X1 U2129 ( .IN1(\U292/DATA1_7 ), .IN2(n14410), .IN3(n14402), .IN4(n9885), .IN5(\U297/DATA1_7 ), .IN6(n14387), .Q(n9884) );
  OR2X1 U2130 ( .IN1(n9886), .IN2(n9887), .Q(n9885) );
  AO221X1 U2131 ( .IN1(\U327/DATA1_7 ), .IN2(n14376), .IN3(\U332/DATA1_7 ), 
        .IN4(n14368), .IN5(n9888), .Q(n9887) );
  AO22X1 U2132 ( .IN1(\U302/DATA1_7 ), .IN2(n14191), .IN3(\U332/DATA2_7 ), 
        .IN4(n14363), .Q(n9888) );
  AO221X1 U2133 ( .IN1(\U307/DATA1_7 ), .IN2(n14354), .IN3(\U322/DATA1_7 ), 
        .IN4(n14338), .IN5(n9889), .Q(n9886) );
  AO22X1 U2134 ( .IN1(\U312/DATA1_7 ), .IN2(n14328), .IN3(\U317/DATA1_7 ), 
        .IN4(n14318), .Q(n9889) );
  AO221X1 U2135 ( .IN1(n5588), .IN2(n14247), .IN3(\U287/DATA1_6 ), .IN4(n14196), .IN5(n9890), .Q(n13262) );
  AO222X1 U2136 ( .IN1(\U292/DATA1_6 ), .IN2(n14410), .IN3(n14402), .IN4(n9891), .IN5(p___constant_11x11xf32_5_8[6]), .IN6(n14388), .Q(n9890) );
  OR2X1 U2137 ( .IN1(n9892), .IN2(n9893), .Q(n9891) );
  AO221X1 U2138 ( .IN1(\U327/DATA1_6 ), .IN2(n14377), .IN3(\U332/DATA1_6 ), 
        .IN4(n14368), .IN5(n9894), .Q(n9893) );
  AO22X1 U2139 ( .IN1(\U302/DATA1_6 ), .IN2(n14191), .IN3(\U332/DATA2_6 ), 
        .IN4(n14355), .Q(n9894) );
  AO221X1 U2140 ( .IN1(\U307/DATA1_6 ), .IN2(n14346), .IN3(\U322/DATA1_6 ), 
        .IN4(n14338), .IN5(n9895), .Q(n9892) );
  AO22X1 U2141 ( .IN1(\U312/DATA1_6 ), .IN2(n14328), .IN3(\U317/DATA1_6 ), 
        .IN4(n14318), .Q(n9895) );
  AO221X1 U2142 ( .IN1(n5587), .IN2(n14247), .IN3(\U287/DATA1_5 ), .IN4(n14196), .IN5(n9896), .Q(n13263) );
  AO222X1 U2143 ( .IN1(\U292/DATA1_5 ), .IN2(n14410), .IN3(n14402), .IN4(n9897), .IN5(p___constant_11x11xf32_5_8[5]), .IN6(n14386), .Q(n9896) );
  OR2X1 U2144 ( .IN1(n9898), .IN2(n9899), .Q(n9897) );
  AO221X1 U2145 ( .IN1(\U327/DATA1_5 ), .IN2(n14383), .IN3(\U332/DATA1_5 ), 
        .IN4(n14368), .IN5(n9900), .Q(n9899) );
  AO22X1 U2146 ( .IN1(\U302/DATA1_5 ), .IN2(n14190), .IN3(\U332/DATA2_5 ), 
        .IN4(n14360), .Q(n9900) );
  AO221X1 U2147 ( .IN1(\U307/DATA1_5 ), .IN2(n14347), .IN3(\U322/DATA1_5 ), 
        .IN4(n14338), .IN5(n9901), .Q(n9898) );
  AO22X1 U2148 ( .IN1(\U312/DATA1_5 ), .IN2(n14328), .IN3(\U317/DATA1_5 ), 
        .IN4(n14318), .Q(n9901) );
  AO221X1 U2149 ( .IN1(n5586), .IN2(n14247), .IN3(\U287/DATA1_4 ), .IN4(n14196), .IN5(n9902), .Q(n13264) );
  AO222X1 U2150 ( .IN1(\U292/DATA1_4 ), .IN2(n14410), .IN3(n14402), .IN4(n9903), .IN5(p___constant_11x11xf32_5_8[4]), .IN6(n14394), .Q(n9902) );
  OR2X1 U2151 ( .IN1(n9904), .IN2(n9905), .Q(n9903) );
  AO221X1 U2152 ( .IN1(\U327/DATA1_4 ), .IN2(n14378), .IN3(\U332/DATA1_4 ), 
        .IN4(n14368), .IN5(n9906), .Q(n9905) );
  AO22X1 U2153 ( .IN1(\U302/DATA1_4 ), .IN2(n14192), .IN3(\U332/DATA2_4 ), 
        .IN4(n14357), .Q(n9906) );
  AO221X1 U2154 ( .IN1(p___constant_11x11xf32_5_6[4]), .IN2(n14345), .IN3(
        \U322/DATA1_4 ), .IN4(n14338), .IN5(n9907), .Q(n9904) );
  AO22X1 U2155 ( .IN1(\U312/DATA1_4 ), .IN2(n14328), .IN3(\U317/DATA1_4 ), 
        .IN4(n14318), .Q(n9907) );
  AO221X1 U2156 ( .IN1(n5585), .IN2(n14247), .IN3(\U287/DATA1_3 ), .IN4(n14196), .IN5(n9908), .Q(n13265) );
  AO222X1 U2157 ( .IN1(\U292/DATA1_3 ), .IN2(n14410), .IN3(n14402), .IN4(n9909), .IN5(p___constant_11x11xf32_5_8[3]), .IN6(n14389), .Q(n9908) );
  OR2X1 U2158 ( .IN1(n9910), .IN2(n9911), .Q(n9909) );
  AO221X1 U2159 ( .IN1(\U327/DATA1_3 ), .IN2(n14384), .IN3(\U332/DATA1_3 ), 
        .IN4(n14368), .IN5(n9912), .Q(n9911) );
  AO22X1 U2160 ( .IN1(\U302/DATA1_3 ), .IN2(n14186), .IN3(\U332/DATA2_3 ), 
        .IN4(n14363), .Q(n9912) );
  AO221X1 U2161 ( .IN1(p___constant_11x11xf32_5_6[3]), .IN2(n14348), .IN3(
        \U322/DATA1_3 ), .IN4(n14338), .IN5(n9913), .Q(n9910) );
  AO22X1 U2162 ( .IN1(\U312/DATA1_3 ), .IN2(n14328), .IN3(\U317/DATA1_3 ), 
        .IN4(n14318), .Q(n9913) );
  AO221X1 U2163 ( .IN1(n5584), .IN2(n14247), .IN3(\U287/DATA1_2 ), .IN4(n14196), .IN5(n9914), .Q(n13266) );
  AO222X1 U2164 ( .IN1(\U292/DATA1_2 ), .IN2(n14410), .IN3(n14402), .IN4(n9915), .IN5(p___constant_11x11xf32_5_8[2]), .IN6(n14394), .Q(n9914) );
  OR2X1 U2165 ( .IN1(n9916), .IN2(n9917), .Q(n9915) );
  AO221X1 U2166 ( .IN1(\U327/DATA1_2 ), .IN2(n14385), .IN3(\U332/DATA1_2 ), 
        .IN4(n14368), .IN5(n9918), .Q(n9917) );
  AO22X1 U2167 ( .IN1(\U302/DATA1_2 ), .IN2(n14257), .IN3(\U332/DATA2_2 ), 
        .IN4(n14361), .Q(n9918) );
  AO221X1 U2168 ( .IN1(p___constant_11x11xf32_5_6[2]), .IN2(n14349), .IN3(
        p___constant_11x11xf32_5_3[2]), .IN4(n14338), .IN5(n9919), .Q(n9916)
         );
  AO22X1 U2169 ( .IN1(\U312/DATA1_2 ), .IN2(n14328), .IN3(\U317/DATA1_2 ), 
        .IN4(n14318), .Q(n9919) );
  AO221X1 U2170 ( .IN1(n5583), .IN2(n14246), .IN3(
        p___constant_11x11xf32_5_10[1]), .IN4(n14196), .IN5(n9920), .Q(n13267)
         );
  AO222X1 U2171 ( .IN1(\U292/DATA1_1 ), .IN2(n14410), .IN3(n14402), .IN4(n9921), .IN5(p___constant_11x11xf32_5_8[1]), .IN6(n14388), .Q(n9920) );
  OR2X1 U2172 ( .IN1(n9922), .IN2(n9923), .Q(n9921) );
  AO221X1 U2173 ( .IN1(p___constant_11x11xf32_5_2[1]), .IN2(n14377), .IN3(
        \U332/DATA1_1 ), .IN4(n14368), .IN5(n9924), .Q(n9923) );
  AO22X1 U2174 ( .IN1(\U302/DATA1_1 ), .IN2(n14189), .IN3(\U332/DATA2_1 ), 
        .IN4(n14357), .Q(n9924) );
  AO221X1 U2175 ( .IN1(p___constant_11x11xf32_5_6[1]), .IN2(n14346), .IN3(
        p___constant_11x11xf32_5_3[1]), .IN4(n14338), .IN5(n9925), .Q(n9922)
         );
  AO22X1 U2176 ( .IN1(\U312/DATA1_1 ), .IN2(n14328), .IN3(\U317/DATA1_1 ), 
        .IN4(n14318), .Q(n9925) );
  AO221X1 U2177 ( .IN1(n5582), .IN2(n14250), .IN3(
        p___constant_11x11xf32_5_10[0]), .IN4(n14196), .IN5(n9926), .Q(n13268)
         );
  AO222X1 U2178 ( .IN1(p___constant_11x11xf32_5_9[0]), .IN2(n14410), .IN3(
        n14402), .IN4(n9927), .IN5(p___constant_11x11xf32_5_8[0]), .IN6(n14390), .Q(n9926) );
  OR2X1 U2179 ( .IN1(n9928), .IN2(n9929), .Q(n9927) );
  AO221X1 U2180 ( .IN1(p___constant_11x11xf32_5_2[0]), .IN2(n14379), .IN3(
        p___constant_11x11xf32_5_1[0]), .IN4(n14368), .IN5(n9930), .Q(n9929)
         );
  AO22X1 U2181 ( .IN1(p___constant_11x11xf32_5_7[0]), .IN2(n14256), .IN3(
        p___constant_11x11xf32_5_0[0]), .IN4(n14357), .Q(n9930) );
  AO221X1 U2182 ( .IN1(p___constant_11x11xf32_5_6[0]), .IN2(n14352), .IN3(
        p___constant_11x11xf32_5_3[0]), .IN4(n14338), .IN5(n9931), .Q(n9928)
         );
  AO22X1 U2183 ( .IN1(p___constant_11x11xf32_5_5[0]), .IN2(n14328), .IN3(
        p___constant_11x11xf32_5_4[0]), .IN4(n14318), .Q(n9931) );
  AO21X1 U2184 ( .IN1(n14239), .IN2(n13760), .IN3(n9529), .Q(n13269) );
  AO21X1 U2185 ( .IN1(n14239), .IN2(n13613), .IN3(n9531), .Q(n13270) );
  AO21X1 U2186 ( .IN1(n14240), .IN2(n14072), .IN3(n9533), .Q(n13271) );
  AO21X1 U2188 ( .IN1(n5602), .IN2(n14241), .IN3(n9534), .Q(n13272) );
  AO21X1 U2189 ( .IN1(n5601), .IN2(n14241), .IN3(n9535), .Q(n13273) );
  AO21X1 U2190 ( .IN1(n5600), .IN2(n14242), .IN3(n9536), .Q(n13274) );
  AO21X1 U2191 ( .IN1(n5599), .IN2(n14246), .IN3(n9537), .Q(n13275) );
  AO21X1 U2192 ( .IN1(n5598), .IN2(n14246), .IN3(n9538), .Q(n13276) );
  AO21X1 U2193 ( .IN1(n5597), .IN2(n14246), .IN3(n9540), .Q(n13277) );
  AO21X1 U2194 ( .IN1(n5596), .IN2(n14246), .IN3(n9542), .Q(n13278) );
  AO21X1 U2195 ( .IN1(n5595), .IN2(n14246), .IN3(n9544), .Q(n13279) );
  AO221X1 U2197 ( .IN1(n14237), .IN2(n13912), .IN3(\U346/DATA1_11 ), .IN4(
        n14197), .IN5(n9936), .Q(n13281) );
  AO222X1 U2198 ( .IN1(\U351/DATA1_11 ), .IN2(n14410), .IN3(n14403), .IN4(
        n9937), .IN5(\U356/DATA1_11 ), .IN6(n14390), .Q(n9936) );
  OR2X1 U2199 ( .IN1(n9938), .IN2(n9939), .Q(n9937) );
  AO221X1 U2200 ( .IN1(\U386/DATA1_11 ), .IN2(n14380), .IN3(\U391/DATA1_11 ), 
        .IN4(n14367), .IN5(n9940), .Q(n9939) );
  AO22X1 U2201 ( .IN1(\U361/DATA1_11 ), .IN2(n14255), .IN3(\U391/DATA2_11 ), 
        .IN4(n14357), .Q(n9940) );
  AO221X1 U2202 ( .IN1(\U366/DATA1_11 ), .IN2(n14349), .IN3(\U381/DATA1_11 ), 
        .IN4(n14337), .IN5(n9941), .Q(n9938) );
  AO22X1 U2203 ( .IN1(\U371/DATA1_11 ), .IN2(n14327), .IN3(\U376/DATA1_11 ), 
        .IN4(n14317), .Q(n9941) );
  AO221X1 U2205 ( .IN1(n14237), .IN2(n13902), .IN3(\U346/DATA1_10 ), .IN4(
        n14197), .IN5(n9943), .Q(n13282) );
  AO222X1 U2206 ( .IN1(\U351/DATA1_10 ), .IN2(n14410), .IN3(n14403), .IN4(
        n9944), .IN5(\U356/DATA1_10 ), .IN6(n14390), .Q(n9943) );
  OR2X1 U2207 ( .IN1(n9945), .IN2(n9946), .Q(n9944) );
  AO221X1 U2208 ( .IN1(\U386/DATA1_10 ), .IN2(n14380), .IN3(\U391/DATA1_10 ), 
        .IN4(n14367), .IN5(n9947), .Q(n9946) );
  AO22X1 U2209 ( .IN1(\U361/DATA1_10 ), .IN2(n14186), .IN3(\U391/DATA2_10 ), 
        .IN4(n14357), .Q(n9947) );
  AO221X1 U2210 ( .IN1(\U366/DATA1_10 ), .IN2(n14349), .IN3(\U381/DATA1_10 ), 
        .IN4(n14337), .IN5(n9948), .Q(n9945) );
  AO22X1 U2211 ( .IN1(\U371/DATA1_10 ), .IN2(n14327), .IN3(\U376/DATA1_10 ), 
        .IN4(n14317), .Q(n9948) );
  AO221X1 U2212 ( .IN1(n14237), .IN2(n14044), .IN3(\U346/DATA1_9 ), .IN4(
        n14197), .IN5(n9950), .Q(n13283) );
  AO222X1 U2213 ( .IN1(\U351/DATA1_9 ), .IN2(n14410), .IN3(n14403), .IN4(n9951), .IN5(\U356/DATA1_9 ), .IN6(n14390), .Q(n9950) );
  OR2X1 U2214 ( .IN1(n9952), .IN2(n9953), .Q(n9951) );
  AO221X1 U2215 ( .IN1(\U386/DATA1_9 ), .IN2(n14380), .IN3(\U391/DATA1_9 ), 
        .IN4(n14367), .IN5(n9954), .Q(n9953) );
  AO22X1 U2216 ( .IN1(\U361/DATA1_9 ), .IN2(n14190), .IN3(\U391/DATA2_9 ), 
        .IN4(n14357), .Q(n9954) );
  AO221X1 U2217 ( .IN1(\U366/DATA1_9 ), .IN2(n14349), .IN3(\U381/DATA1_9 ), 
        .IN4(n14337), .IN5(n9955), .Q(n9952) );
  AO22X1 U2218 ( .IN1(\U371/DATA1_9 ), .IN2(n14327), .IN3(\U376/DATA1_9 ), 
        .IN4(n14317), .Q(n9955) );
  AO221X1 U2220 ( .IN1(n5662), .IN2(n14249), .IN3(\U346/DATA1_8 ), .IN4(n14197), .IN5(n9956), .Q(n13284) );
  AO222X1 U2221 ( .IN1(\U351/DATA1_8 ), .IN2(n14411), .IN3(n14403), .IN4(n9957), .IN5(\U356/DATA1_8 ), .IN6(n14390), .Q(n9956) );
  OR2X1 U2222 ( .IN1(n9958), .IN2(n9959), .Q(n9957) );
  AO221X1 U2223 ( .IN1(\U386/DATA1_8 ), .IN2(n14380), .IN3(\U391/DATA1_8 ), 
        .IN4(n14367), .IN5(n9960), .Q(n9959) );
  AO22X1 U2224 ( .IN1(\U361/DATA1_8 ), .IN2(n14193), .IN3(\U391/DATA2_8 ), 
        .IN4(n14357), .Q(n9960) );
  AO221X1 U2225 ( .IN1(\U366/DATA1_8 ), .IN2(n14349), .IN3(\U381/DATA1_8 ), 
        .IN4(n14337), .IN5(n9961), .Q(n9958) );
  AO22X1 U2226 ( .IN1(\U371/DATA1_8 ), .IN2(n14327), .IN3(\U376/DATA1_8 ), 
        .IN4(n14317), .Q(n9961) );
  AO221X1 U2227 ( .IN1(n5661), .IN2(n14248), .IN3(\U346/DATA1_7 ), .IN4(n14197), .IN5(n9962), .Q(n13285) );
  AO222X1 U2228 ( .IN1(\U351/DATA1_7 ), .IN2(n14411), .IN3(n14403), .IN4(n9963), .IN5(\U356/DATA1_7 ), .IN6(n14390), .Q(n9962) );
  OR2X1 U2229 ( .IN1(n9964), .IN2(n9965), .Q(n9963) );
  AO221X1 U2230 ( .IN1(\U386/DATA1_7 ), .IN2(n14380), .IN3(\U391/DATA1_7 ), 
        .IN4(n14367), .IN5(n9966), .Q(n9965) );
  AO22X1 U2231 ( .IN1(\U361/DATA1_7 ), .IN2(n14257), .IN3(\U391/DATA2_7 ), 
        .IN4(n14357), .Q(n9966) );
  AO221X1 U2232 ( .IN1(\U366/DATA1_7 ), .IN2(n14349), .IN3(\U381/DATA1_7 ), 
        .IN4(n14337), .IN5(n9967), .Q(n9964) );
  AO22X1 U2233 ( .IN1(\U371/DATA1_7 ), .IN2(n14327), .IN3(\U376/DATA1_7 ), 
        .IN4(n14317), .Q(n9967) );
  AO221X1 U2234 ( .IN1(n5660), .IN2(n14248), .IN3(\U346/DATA1_6 ), .IN4(n14197), .IN5(n9968), .Q(n13286) );
  AO222X1 U2235 ( .IN1(\U351/DATA1_6 ), .IN2(n14411), .IN3(n14403), .IN4(n9969), .IN5(\U356/DATA1_6 ), .IN6(n14390), .Q(n9968) );
  OR2X1 U2236 ( .IN1(n9970), .IN2(n9971), .Q(n9969) );
  AO221X1 U2237 ( .IN1(\U386/DATA1_6 ), .IN2(n14380), .IN3(\U391/DATA1_6 ), 
        .IN4(n14367), .IN5(n9972), .Q(n9971) );
  AO22X1 U2238 ( .IN1(\U361/DATA1_6 ), .IN2(n14189), .IN3(\U391/DATA2_6 ), 
        .IN4(n14357), .Q(n9972) );
  AO221X1 U2239 ( .IN1(\U366/DATA1_6 ), .IN2(n14349), .IN3(\U381/DATA1_6 ), 
        .IN4(n14337), .IN5(n9973), .Q(n9970) );
  AO22X1 U2240 ( .IN1(\U371/DATA1_6 ), .IN2(n14327), .IN3(\U376/DATA1_6 ), 
        .IN4(n14317), .Q(n9973) );
  AO221X1 U2241 ( .IN1(n5659), .IN2(n14248), .IN3(\U346/DATA1_5 ), .IN4(n14197), .IN5(n9974), .Q(n13287) );
  AO222X1 U2242 ( .IN1(\U351/DATA1_5 ), .IN2(n14411), .IN3(n14403), .IN4(n9975), .IN5(\U356/DATA1_5 ), .IN6(n14390), .Q(n9974) );
  OR2X1 U2243 ( .IN1(n9976), .IN2(n9977), .Q(n9975) );
  AO221X1 U2244 ( .IN1(\U386/DATA1_5 ), .IN2(n14380), .IN3(\U391/DATA1_5 ), 
        .IN4(n14367), .IN5(n9978), .Q(n9977) );
  AO22X1 U2245 ( .IN1(\U361/DATA1_5 ), .IN2(n14192), .IN3(\U391/DATA2_5 ), 
        .IN4(n14357), .Q(n9978) );
  AO221X1 U2246 ( .IN1(\U366/DATA1_5 ), .IN2(n14349), .IN3(\U381/DATA1_5 ), 
        .IN4(n14337), .IN5(n9979), .Q(n9976) );
  AO22X1 U2247 ( .IN1(\U371/DATA1_5 ), .IN2(n14327), .IN3(\U376/DATA1_5 ), 
        .IN4(n14317), .Q(n9979) );
  AO221X1 U2248 ( .IN1(n5658), .IN2(n14249), .IN3(
        p___constant_11x11xf32_4_10[4]), .IN4(n14197), .IN5(n9980), .Q(n13288)
         );
  AO222X1 U2249 ( .IN1(\U351/DATA1_4 ), .IN2(n14411), .IN3(n14403), .IN4(n9981), .IN5(\U356/DATA1_4 ), .IN6(n14390), .Q(n9980) );
  OR2X1 U2250 ( .IN1(n9982), .IN2(n9983), .Q(n9981) );
  AO221X1 U2251 ( .IN1(\U386/DATA1_4 ), .IN2(n14380), .IN3(\U391/DATA1_4 ), 
        .IN4(n14367), .IN5(n9984), .Q(n9983) );
  AO22X1 U2252 ( .IN1(\U361/DATA1_4 ), .IN2(n14254), .IN3(\U391/DATA2_4 ), 
        .IN4(n14357), .Q(n9984) );
  AO221X1 U2253 ( .IN1(\U366/DATA1_4 ), .IN2(n14349), .IN3(\U381/DATA1_4 ), 
        .IN4(n14337), .IN5(n9985), .Q(n9982) );
  AO22X1 U2254 ( .IN1(\U371/DATA1_4 ), .IN2(n14327), .IN3(\U376/DATA1_4 ), 
        .IN4(n14317), .Q(n9985) );
  AO221X1 U2255 ( .IN1(n5657), .IN2(n14249), .IN3(
        p___constant_11x11xf32_4_10[3]), .IN4(n14197), .IN5(n9986), .Q(n13289)
         );
  AO222X1 U2256 ( .IN1(\U351/DATA1_3 ), .IN2(n14411), .IN3(n14403), .IN4(n9987), .IN5(\U356/DATA1_3 ), .IN6(n14390), .Q(n9986) );
  OR2X1 U2257 ( .IN1(n9988), .IN2(n9989), .Q(n9987) );
  AO221X1 U2258 ( .IN1(\U386/DATA1_3 ), .IN2(n14380), .IN3(\U391/DATA1_3 ), 
        .IN4(n14367), .IN5(n9990), .Q(n9989) );
  AO22X1 U2259 ( .IN1(\U361/DATA1_3 ), .IN2(n14190), .IN3(\U391/DATA2_3 ), 
        .IN4(n14357), .Q(n9990) );
  AO221X1 U2260 ( .IN1(\U366/DATA1_3 ), .IN2(n14349), .IN3(\U381/DATA1_3 ), 
        .IN4(n14337), .IN5(n9991), .Q(n9988) );
  AO22X1 U2261 ( .IN1(\U371/DATA1_3 ), .IN2(n14327), .IN3(\U376/DATA1_3 ), 
        .IN4(n14317), .Q(n9991) );
  AO221X1 U2262 ( .IN1(n5656), .IN2(n14249), .IN3(
        p___constant_11x11xf32_4_10[2]), .IN4(n14197), .IN5(n9992), .Q(n13290)
         );
  AO222X1 U2263 ( .IN1(\U351/DATA1_2 ), .IN2(n14411), .IN3(n14403), .IN4(n9993), .IN5(\U356/DATA1_2 ), .IN6(n14390), .Q(n9992) );
  OR2X1 U2264 ( .IN1(n9994), .IN2(n9995), .Q(n9993) );
  AO221X1 U2265 ( .IN1(\U386/DATA1_2 ), .IN2(n14380), .IN3(\U391/DATA1_2 ), 
        .IN4(n14367), .IN5(n9996), .Q(n9995) );
  AO22X1 U2266 ( .IN1(p___constant_11x11xf32_4_7[2]), .IN2(n14191), .IN3(
        \U391/DATA2_2 ), .IN4(n14357), .Q(n9996) );
  AO221X1 U2267 ( .IN1(\U366/DATA1_2 ), .IN2(n14349), .IN3(\U381/DATA1_2 ), 
        .IN4(n14337), .IN5(n9997), .Q(n9994) );
  AO22X1 U2268 ( .IN1(\U371/DATA1_2 ), .IN2(n14327), .IN3(\U376/DATA1_2 ), 
        .IN4(n14317), .Q(n9997) );
  AO221X1 U2269 ( .IN1(n5655), .IN2(n14249), .IN3(
        p___constant_11x11xf32_4_10[1]), .IN4(n14197), .IN5(n9998), .Q(n13291)
         );
  AO222X1 U2270 ( .IN1(\U351/DATA1_1 ), .IN2(n14411), .IN3(n14403), .IN4(n9999), .IN5(\U356/DATA1_1 ), .IN6(n14390), .Q(n9998) );
  OR2X1 U2271 ( .IN1(n10000), .IN2(n10001), .Q(n9999) );
  AO221X1 U2272 ( .IN1(\U386/DATA1_1 ), .IN2(n14380), .IN3(\U391/DATA1_1 ), 
        .IN4(n14367), .IN5(n10002), .Q(n10001) );
  AO22X1 U2273 ( .IN1(p___constant_11x11xf32_4_7[1]), .IN2(n14190), .IN3(
        \U391/DATA2_1 ), .IN4(n14357), .Q(n10002) );
  AO221X1 U2274 ( .IN1(\U366/DATA1_1 ), .IN2(n14349), .IN3(\U381/DATA1_1 ), 
        .IN4(n14337), .IN5(n10003), .Q(n10000) );
  AO22X1 U2275 ( .IN1(\U371/DATA1_1 ), .IN2(n14327), .IN3(\U376/DATA1_1 ), 
        .IN4(n14317), .Q(n10003) );
  AO221X1 U2276 ( .IN1(n5654), .IN2(n14249), .IN3(
        p___constant_11x11xf32_4_10[0]), .IN4(n13736), .IN5(n10004), .Q(n13292) );
  AO222X1 U2277 ( .IN1(p___constant_11x11xf32_4_9[0]), .IN2(n14411), .IN3(
        n14403), .IN4(n10005), .IN5(p___constant_11x11xf32_4_8[0]), .IN6(
        n14390), .Q(n10004) );
  OR2X1 U2278 ( .IN1(n10006), .IN2(n10007), .Q(n10005) );
  AO221X1 U2279 ( .IN1(\U386/DATA1_0 ), .IN2(n14380), .IN3(\U391/DATA1_0 ), 
        .IN4(n14367), .IN5(n10008), .Q(n10007) );
  AO22X1 U2280 ( .IN1(p___constant_11x11xf32_4_7[0]), .IN2(n14254), .IN3(
        \U391/DATA2_0 ), .IN4(n14357), .Q(n10008) );
  AO221X1 U2281 ( .IN1(\U366/DATA1_0 ), .IN2(n14349), .IN3(\U381/DATA1_0 ), 
        .IN4(n14337), .IN5(n10009), .Q(n10006) );
  AO22X1 U2282 ( .IN1(\U371/DATA1_0 ), .IN2(n14327), .IN3(\U376/DATA1_0 ), 
        .IN4(n14317), .Q(n10009) );
  AO21X1 U2283 ( .IN1(n14240), .IN2(n13759), .IN3(n9529), .Q(n13293) );
  AO21X1 U2284 ( .IN1(n14240), .IN2(n13612), .IN3(n9531), .Q(n13294) );
  AO21X1 U2285 ( .IN1(n14241), .IN2(n14071), .IN3(n9533), .Q(n13295) );
  AO21X1 U2287 ( .IN1(n5674), .IN2(n14905), .IN3(n9534), .Q(n13296) );
  AO21X1 U2288 ( .IN1(n5673), .IN2(n14246), .IN3(n9535), .Q(n13297) );
  AO21X1 U2289 ( .IN1(n5672), .IN2(n14246), .IN3(n9536), .Q(n13298) );
  AO21X1 U2290 ( .IN1(n5671), .IN2(n14246), .IN3(n9537), .Q(n13299) );
  AO21X1 U2291 ( .IN1(n5670), .IN2(n14246), .IN3(n9538), .Q(n13300) );
  AO21X1 U2292 ( .IN1(n5669), .IN2(n14246), .IN3(n9540), .Q(n13301) );
  AO21X1 U2293 ( .IN1(n5668), .IN2(n14246), .IN3(n9542), .Q(n13302) );
  AO21X1 U2294 ( .IN1(n5667), .IN2(n14246), .IN3(n9544), .Q(n13303) );
  AO221X1 U2296 ( .IN1(n14238), .IN2(n13911), .IN3(\U399/DATA1_11 ), .IN4(
        n13736), .IN5(n10014), .Q(n13305) );
  AO222X1 U2297 ( .IN1(\U404/DATA1_11 ), .IN2(n14411), .IN3(n14404), .IN4(
        n10015), .IN5(\U409/DATA1_11 ), .IN6(n14391), .Q(n10014) );
  OR2X1 U2298 ( .IN1(n10016), .IN2(n10017), .Q(n10015) );
  AO221X1 U2299 ( .IN1(\U439/DATA1_11 ), .IN2(n14379), .IN3(\U444/DATA1_11 ), 
        .IN4(n14366), .IN5(n10018), .Q(n10017) );
  AO22X1 U2300 ( .IN1(\U414/DATA1_11 ), .IN2(n14914), .IN3(\U444/DATA2_11 ), 
        .IN4(n14357), .Q(n10018) );
  AO221X1 U2301 ( .IN1(\U419/DATA1_11 ), .IN2(n14348), .IN3(\U434/DATA1_11 ), 
        .IN4(n14336), .IN5(n10019), .Q(n10016) );
  AO22X1 U2302 ( .IN1(\U424/DATA1_11 ), .IN2(n14327), .IN3(\U429/DATA1_11 ), 
        .IN4(n14316), .Q(n10019) );
  AO221X1 U2304 ( .IN1(n14238), .IN2(n13901), .IN3(\U399/DATA1_10 ), .IN4(
        n13736), .IN5(n10021), .Q(n13306) );
  AO222X1 U2305 ( .IN1(\U404/DATA1_10 ), .IN2(n14411), .IN3(n14404), .IN4(
        n10022), .IN5(\U409/DATA1_10 ), .IN6(n14391), .Q(n10021) );
  OR2X1 U2306 ( .IN1(n10023), .IN2(n10024), .Q(n10022) );
  AO221X1 U2307 ( .IN1(\U439/DATA1_10 ), .IN2(n14379), .IN3(\U444/DATA1_10 ), 
        .IN4(n14366), .IN5(n10025), .Q(n10024) );
  AO22X1 U2308 ( .IN1(\U414/DATA1_10 ), .IN2(n14189), .IN3(\U444/DATA2_10 ), 
        .IN4(n14357), .Q(n10025) );
  AO221X1 U2309 ( .IN1(\U419/DATA1_10 ), .IN2(n14348), .IN3(\U434/DATA1_10 ), 
        .IN4(n14336), .IN5(n10026), .Q(n10023) );
  AO22X1 U2310 ( .IN1(\U424/DATA1_10 ), .IN2(n14325), .IN3(\U429/DATA1_10 ), 
        .IN4(n14316), .Q(n10026) );
  AO221X1 U2311 ( .IN1(n14236), .IN2(n14043), .IN3(\U399/DATA1_9 ), .IN4(
        n13736), .IN5(n10028), .Q(n13307) );
  AO222X1 U2312 ( .IN1(\U404/DATA1_9 ), .IN2(n14411), .IN3(n14404), .IN4(
        n10029), .IN5(\U409/DATA1_9 ), .IN6(n14391), .Q(n10028) );
  OR2X1 U2313 ( .IN1(n10030), .IN2(n10031), .Q(n10029) );
  AO221X1 U2314 ( .IN1(\U439/DATA1_9 ), .IN2(n14379), .IN3(\U444/DATA1_9 ), 
        .IN4(n14366), .IN5(n10032), .Q(n10031) );
  AO22X1 U2315 ( .IN1(\U414/DATA1_9 ), .IN2(n14914), .IN3(\U444/DATA2_9 ), 
        .IN4(n14358), .Q(n10032) );
  AO221X1 U2316 ( .IN1(\U419/DATA1_9 ), .IN2(n14348), .IN3(\U434/DATA1_9 ), 
        .IN4(n14336), .IN5(n10033), .Q(n10030) );
  AO22X1 U2317 ( .IN1(\U424/DATA1_9 ), .IN2(n14325), .IN3(\U429/DATA1_9 ), 
        .IN4(n14316), .Q(n10033) );
  AO221X1 U2319 ( .IN1(n5734), .IN2(n14234), .IN3(\U399/DATA1_8 ), .IN4(n13736), .IN5(n10034), .Q(n13308) );
  AO222X1 U2320 ( .IN1(\U404/DATA1_8 ), .IN2(n14411), .IN3(n14404), .IN4(
        n10035), .IN5(\U409/DATA1_8 ), .IN6(n14391), .Q(n10034) );
  OR2X1 U2321 ( .IN1(n10036), .IN2(n10037), .Q(n10035) );
  AO221X1 U2322 ( .IN1(\U439/DATA1_8 ), .IN2(n14379), .IN3(\U444/DATA1_8 ), 
        .IN4(n14366), .IN5(n10038), .Q(n10037) );
  AO22X1 U2323 ( .IN1(\U414/DATA1_8 ), .IN2(n14191), .IN3(\U444/DATA2_8 ), 
        .IN4(n14356), .Q(n10038) );
  AO221X1 U2324 ( .IN1(\U419/DATA1_8 ), .IN2(n14348), .IN3(\U434/DATA1_8 ), 
        .IN4(n14336), .IN5(n10039), .Q(n10036) );
  AO22X1 U2325 ( .IN1(\U424/DATA1_8 ), .IN2(n14326), .IN3(\U429/DATA1_8 ), 
        .IN4(n14316), .Q(n10039) );
  AO221X1 U2326 ( .IN1(n5733), .IN2(n14234), .IN3(\U399/DATA1_7 ), .IN4(n13736), .IN5(n10040), .Q(n13309) );
  AO222X1 U2327 ( .IN1(\U404/DATA1_7 ), .IN2(n14411), .IN3(n14404), .IN4(
        n10041), .IN5(\U409/DATA1_7 ), .IN6(n14391), .Q(n10040) );
  OR2X1 U2328 ( .IN1(n10042), .IN2(n10043), .Q(n10041) );
  AO221X1 U2329 ( .IN1(\U439/DATA1_7 ), .IN2(n14379), .IN3(\U444/DATA1_7 ), 
        .IN4(n14366), .IN5(n10044), .Q(n10043) );
  AO22X1 U2330 ( .IN1(\U414/DATA1_7 ), .IN2(n14191), .IN3(\U444/DATA2_7 ), 
        .IN4(n14361), .Q(n10044) );
  AO221X1 U2331 ( .IN1(\U419/DATA1_7 ), .IN2(n14348), .IN3(\U434/DATA1_7 ), 
        .IN4(n14336), .IN5(n10045), .Q(n10042) );
  AO22X1 U2332 ( .IN1(\U424/DATA1_7 ), .IN2(n14325), .IN3(\U429/DATA1_7 ), 
        .IN4(n14316), .Q(n10045) );
  AO221X1 U2333 ( .IN1(n5732), .IN2(n14905), .IN3(\U399/DATA1_6 ), .IN4(n13736), .IN5(n10046), .Q(n13310) );
  AO222X1 U2334 ( .IN1(\U404/DATA1_6 ), .IN2(n14411), .IN3(n14404), .IN4(
        n10047), .IN5(\U409/DATA1_6 ), .IN6(n14391), .Q(n10046) );
  OR2X1 U2335 ( .IN1(n10048), .IN2(n10049), .Q(n10047) );
  AO221X1 U2336 ( .IN1(\U439/DATA1_6 ), .IN2(n14379), .IN3(\U444/DATA1_6 ), 
        .IN4(n14366), .IN5(n10050), .Q(n10049) );
  AO22X1 U2337 ( .IN1(\U414/DATA1_6 ), .IN2(n14192), .IN3(\U444/DATA2_6 ), 
        .IN4(n14362), .Q(n10050) );
  AO221X1 U2338 ( .IN1(\U419/DATA1_6 ), .IN2(n14348), .IN3(\U434/DATA1_6 ), 
        .IN4(n14336), .IN5(n10051), .Q(n10048) );
  AO22X1 U2339 ( .IN1(\U424/DATA1_6 ), .IN2(n14332), .IN3(\U429/DATA1_6 ), 
        .IN4(n14316), .Q(n10051) );
  AO221X1 U2340 ( .IN1(n5731), .IN2(n14237), .IN3(\U399/DATA1_5 ), .IN4(n14198), .IN5(n10052), .Q(n13311) );
  AO222X1 U2341 ( .IN1(\U404/DATA1_5 ), .IN2(n14412), .IN3(n14404), .IN4(
        n10053), .IN5(\U409/DATA1_5 ), .IN6(n14391), .Q(n10052) );
  OR2X1 U2342 ( .IN1(n10054), .IN2(n10055), .Q(n10053) );
  AO221X1 U2343 ( .IN1(\U439/DATA1_5 ), .IN2(n14379), .IN3(\U444/DATA1_5 ), 
        .IN4(n14366), .IN5(n10056), .Q(n10055) );
  AO22X1 U2344 ( .IN1(\U414/DATA1_5 ), .IN2(n14192), .IN3(\U444/DATA2_5 ), 
        .IN4(n14363), .Q(n10056) );
  AO221X1 U2345 ( .IN1(\U419/DATA1_5 ), .IN2(n14348), .IN3(\U434/DATA1_5 ), 
        .IN4(n14336), .IN5(n10057), .Q(n10054) );
  AO22X1 U2346 ( .IN1(\U424/DATA1_5 ), .IN2(n14333), .IN3(\U429/DATA1_5 ), 
        .IN4(n14316), .Q(n10057) );
  AO221X1 U2347 ( .IN1(n5730), .IN2(n14250), .IN3(\U399/DATA1_4 ), .IN4(n14198), .IN5(n10058), .Q(n13312) );
  AO222X1 U2348 ( .IN1(\U404/DATA1_4 ), .IN2(n14412), .IN3(n14404), .IN4(
        n10059), .IN5(\U409/DATA1_4 ), .IN6(n14391), .Q(n10058) );
  OR2X1 U2349 ( .IN1(n10060), .IN2(n10061), .Q(n10059) );
  AO221X1 U2350 ( .IN1(\U439/DATA1_4 ), .IN2(n14379), .IN3(\U444/DATA1_4 ), 
        .IN4(n14366), .IN5(n10062), .Q(n10061) );
  AO22X1 U2351 ( .IN1(\U414/DATA1_4 ), .IN2(n14191), .IN3(\U444/DATA2_4 ), 
        .IN4(n14363), .Q(n10062) );
  AO221X1 U2352 ( .IN1(\U419/DATA1_4 ), .IN2(n14348), .IN3(\U434/DATA1_4 ), 
        .IN4(n14336), .IN5(n10063), .Q(n10060) );
  AO22X1 U2353 ( .IN1(\U424/DATA1_4 ), .IN2(n14329), .IN3(\U429/DATA1_4 ), 
        .IN4(n14316), .Q(n10063) );
  AO221X1 U2354 ( .IN1(n5729), .IN2(n14241), .IN3(\U399/DATA1_3 ), .IN4(n14198), .IN5(n10064), .Q(n13313) );
  AO222X1 U2355 ( .IN1(\U404/DATA1_3 ), .IN2(n14412), .IN3(n14404), .IN4(
        n10065), .IN5(\U409/DATA1_3 ), .IN6(n14391), .Q(n10064) );
  OR2X1 U2356 ( .IN1(n10066), .IN2(n10067), .Q(n10065) );
  AO221X1 U2357 ( .IN1(\U439/DATA1_3 ), .IN2(n14379), .IN3(\U444/DATA1_3 ), 
        .IN4(n14366), .IN5(n10068), .Q(n10067) );
  AO22X1 U2358 ( .IN1(\U414/DATA1_3 ), .IN2(n14192), .IN3(\U444/DATA2_3 ), 
        .IN4(n14361), .Q(n10068) );
  AO221X1 U2359 ( .IN1(\U419/DATA1_3 ), .IN2(n14348), .IN3(\U434/DATA1_3 ), 
        .IN4(n14336), .IN5(n10069), .Q(n10066) );
  AO22X1 U2360 ( .IN1(\U424/DATA1_3 ), .IN2(n14331), .IN3(\U429/DATA1_3 ), 
        .IN4(n14316), .Q(n10069) );
  AO221X1 U2361 ( .IN1(n5728), .IN2(n14240), .IN3(\U399/DATA1_2 ), .IN4(n14198), .IN5(n10070), .Q(n13314) );
  AO222X1 U2362 ( .IN1(\U404/DATA1_2 ), .IN2(n14412), .IN3(n14404), .IN4(
        n10071), .IN5(\U409/DATA1_2 ), .IN6(n14391), .Q(n10070) );
  OR2X1 U2363 ( .IN1(n10072), .IN2(n10073), .Q(n10071) );
  AO221X1 U2364 ( .IN1(\U439/DATA1_2 ), .IN2(n14379), .IN3(\U444/DATA1_2 ), 
        .IN4(n14366), .IN5(n10074), .Q(n10073) );
  AO22X1 U2365 ( .IN1(\U414/DATA1_2 ), .IN2(n14186), .IN3(\U444/DATA2_2 ), 
        .IN4(n14361), .Q(n10074) );
  AO221X1 U2366 ( .IN1(\U419/DATA1_2 ), .IN2(n14348), .IN3(\U434/DATA1_2 ), 
        .IN4(n14336), .IN5(n10075), .Q(n10072) );
  AO22X1 U2367 ( .IN1(\U424/DATA1_2 ), .IN2(n14325), .IN3(\U429/DATA1_2 ), 
        .IN4(n14316), .Q(n10075) );
  AO221X1 U2368 ( .IN1(n5727), .IN2(n14248), .IN3(\U399/DATA1_1 ), .IN4(n14198), .IN5(n10076), .Q(n13315) );
  AO222X1 U2369 ( .IN1(\U404/DATA1_1 ), .IN2(n14412), .IN3(n14404), .IN4(
        n10077), .IN5(\U409/DATA1_1 ), .IN6(n14391), .Q(n10076) );
  OR2X1 U2370 ( .IN1(n10078), .IN2(n10079), .Q(n10077) );
  AO221X1 U2371 ( .IN1(\U439/DATA1_1 ), .IN2(n14379), .IN3(\U444/DATA1_1 ), 
        .IN4(n14366), .IN5(n10080), .Q(n10079) );
  AO22X1 U2372 ( .IN1(\U414/DATA1_1 ), .IN2(n14914), .IN3(\U444/DATA2_1 ), 
        .IN4(n14359), .Q(n10080) );
  AO221X1 U2373 ( .IN1(\U419/DATA1_1 ), .IN2(n14348), .IN3(\U434/DATA1_1 ), 
        .IN4(n14336), .IN5(n10081), .Q(n10078) );
  AO22X1 U2374 ( .IN1(\U424/DATA1_1 ), .IN2(n14328), .IN3(\U429/DATA1_1 ), 
        .IN4(n14316), .Q(n10081) );
  AO221X1 U2375 ( .IN1(n5726), .IN2(n14237), .IN3(\U399/DATA1_0 ), .IN4(n14198), .IN5(n10082), .Q(n13316) );
  AO222X1 U2376 ( .IN1(\U404/DATA1_0 ), .IN2(n14412), .IN3(n14404), .IN4(
        n10083), .IN5(\U409/DATA1_0 ), .IN6(n14391), .Q(n10082) );
  OR2X1 U2377 ( .IN1(n10084), .IN2(n10085), .Q(n10083) );
  AO221X1 U2378 ( .IN1(\U439/DATA1_0 ), .IN2(n14379), .IN3(\U444/DATA1_0 ), 
        .IN4(n14366), .IN5(n10086), .Q(n10085) );
  AO22X1 U2379 ( .IN1(\U414/DATA1_0 ), .IN2(n14191), .IN3(\U444/DATA2_0 ), 
        .IN4(n14363), .Q(n10086) );
  AO221X1 U2380 ( .IN1(\U419/DATA1_0 ), .IN2(n14348), .IN3(\U434/DATA1_0 ), 
        .IN4(n14336), .IN5(n10087), .Q(n10084) );
  AO22X1 U2381 ( .IN1(\U424/DATA1_0 ), .IN2(n14330), .IN3(\U429/DATA1_0 ), 
        .IN4(n14316), .Q(n10087) );
  AO21X1 U2382 ( .IN1(n14241), .IN2(n13758), .IN3(n9529), .Q(n13317) );
  AO21X1 U2383 ( .IN1(n14241), .IN2(n13611), .IN3(n9531), .Q(n13318) );
  AO21X1 U2384 ( .IN1(n14241), .IN2(n14070), .IN3(n9533), .Q(n13319) );
  AO21X1 U2386 ( .IN1(n5746), .IN2(n14246), .IN3(n9534), .Q(n13320) );
  AO21X1 U2387 ( .IN1(n5745), .IN2(n14237), .IN3(n9535), .Q(n13321) );
  AO21X1 U2388 ( .IN1(n5744), .IN2(n14234), .IN3(n9536), .Q(n13322) );
  AO21X1 U2389 ( .IN1(n5743), .IN2(n14243), .IN3(n9537), .Q(n13323) );
  AO21X1 U2390 ( .IN1(n5742), .IN2(n14246), .IN3(n9538), .Q(n13324) );
  AO21X1 U2391 ( .IN1(n5741), .IN2(n14244), .IN3(n9540), .Q(n13325) );
  AO21X1 U2392 ( .IN1(n5740), .IN2(n14238), .IN3(n9542), .Q(n13326) );
  AO21X1 U2393 ( .IN1(n5739), .IN2(n14245), .IN3(n9544), .Q(n13327) );
  AO221X1 U2395 ( .IN1(n14237), .IN2(n13910), .IN3(\U455/DATA1_11 ), .IN4(
        n14198), .IN5(n10092), .Q(n13329) );
  AO222X1 U2396 ( .IN1(\U460/DATA1_11 ), .IN2(n14412), .IN3(n14405), .IN4(
        n10093), .IN5(\U465/DATA1_11 ), .IN6(n14392), .Q(n10092) );
  OR2X1 U2397 ( .IN1(n10094), .IN2(n10095), .Q(n10093) );
  AO221X1 U2398 ( .IN1(\U495/DATA1_11 ), .IN2(n14378), .IN3(\U500/DATA1_11 ), 
        .IN4(n14365), .IN5(n10096), .Q(n10095) );
  AO22X1 U2399 ( .IN1(\U470/DATA1_11 ), .IN2(n14254), .IN3(\U500/DATA2_11 ), 
        .IN4(n14361), .Q(n10096) );
  AO221X1 U2400 ( .IN1(\U475/DATA1_11 ), .IN2(n14347), .IN3(\U490/DATA1_11 ), 
        .IN4(n14335), .IN5(n10097), .Q(n10094) );
  AO22X1 U2401 ( .IN1(\U480/DATA1_11 ), .IN2(n14332), .IN3(\U485/DATA1_11 ), 
        .IN4(n14315), .Q(n10097) );
  AO221X1 U2403 ( .IN1(n14237), .IN2(n13900), .IN3(\U455/DATA1_10 ), .IN4(
        n14198), .IN5(n10099), .Q(n13330) );
  AO222X1 U2404 ( .IN1(\U460/DATA1_10 ), .IN2(n14412), .IN3(n14405), .IN4(
        n10100), .IN5(\U465/DATA1_10 ), .IN6(n14392), .Q(n10099) );
  OR2X1 U2405 ( .IN1(n10101), .IN2(n10102), .Q(n10100) );
  AO221X1 U2406 ( .IN1(\U495/DATA1_10 ), .IN2(n14378), .IN3(\U500/DATA1_10 ), 
        .IN4(n14364), .IN5(n10103), .Q(n10102) );
  AO22X1 U2407 ( .IN1(\U470/DATA1_10 ), .IN2(n14190), .IN3(\U500/DATA2_10 ), 
        .IN4(n14362), .Q(n10103) );
  AO221X1 U2408 ( .IN1(\U475/DATA1_10 ), .IN2(n14347), .IN3(\U490/DATA1_10 ), 
        .IN4(n14335), .IN5(n10104), .Q(n10101) );
  AO22X1 U2409 ( .IN1(\U480/DATA1_10 ), .IN2(n14333), .IN3(\U485/DATA1_10 ), 
        .IN4(n14315), .Q(n10104) );
  AO221X1 U2410 ( .IN1(n14236), .IN2(n14042), .IN3(\U455/DATA1_9 ), .IN4(
        n14198), .IN5(n10106), .Q(n13331) );
  AO222X1 U2411 ( .IN1(\U460/DATA1_9 ), .IN2(n14412), .IN3(n14405), .IN4(
        n10107), .IN5(\U465/DATA1_9 ), .IN6(n14392), .Q(n10106) );
  OR2X1 U2412 ( .IN1(n10108), .IN2(n10109), .Q(n10107) );
  AO221X1 U2413 ( .IN1(\U495/DATA1_9 ), .IN2(n14378), .IN3(\U500/DATA1_9 ), 
        .IN4(n14371), .IN5(n10110), .Q(n10109) );
  AO22X1 U2414 ( .IN1(\U470/DATA1_9 ), .IN2(n14257), .IN3(\U500/DATA2_9 ), 
        .IN4(n14360), .Q(n10110) );
  AO221X1 U2415 ( .IN1(\U475/DATA1_9 ), .IN2(n14347), .IN3(\U490/DATA1_9 ), 
        .IN4(n14335), .IN5(n10111), .Q(n10108) );
  AO22X1 U2416 ( .IN1(\U480/DATA1_9 ), .IN2(n14326), .IN3(\U485/DATA1_9 ), 
        .IN4(n14315), .Q(n10111) );
  AO221X1 U2418 ( .IN1(n5806), .IN2(n14239), .IN3(\U455/DATA1_8 ), .IN4(n14198), .IN5(n10112), .Q(n13332) );
  AO222X1 U2419 ( .IN1(\U460/DATA1_8 ), .IN2(n14412), .IN3(n14405), .IN4(
        n10113), .IN5(\U465/DATA1_8 ), .IN6(n14392), .Q(n10112) );
  OR2X1 U2420 ( .IN1(n10114), .IN2(n10115), .Q(n10113) );
  AO221X1 U2421 ( .IN1(\U495/DATA1_8 ), .IN2(n14378), .IN3(\U500/DATA1_8 ), 
        .IN4(n14373), .IN5(n10116), .Q(n10115) );
  AO22X1 U2422 ( .IN1(\U470/DATA1_8 ), .IN2(n14193), .IN3(\U500/DATA2_8 ), 
        .IN4(n14362), .Q(n10116) );
  AO221X1 U2423 ( .IN1(\U475/DATA1_8 ), .IN2(n14347), .IN3(\U490/DATA1_8 ), 
        .IN4(n14335), .IN5(n10117), .Q(n10114) );
  AO22X1 U2424 ( .IN1(\U480/DATA1_8 ), .IN2(n14330), .IN3(\U485/DATA1_8 ), 
        .IN4(n14315), .Q(n10117) );
  AO221X1 U2425 ( .IN1(n5805), .IN2(n14246), .IN3(\U455/DATA1_7 ), .IN4(n14198), .IN5(n10118), .Q(n13333) );
  AO222X1 U2426 ( .IN1(\U460/DATA1_7 ), .IN2(n14412), .IN3(n14405), .IN4(
        n10119), .IN5(\U465/DATA1_7 ), .IN6(n14392), .Q(n10118) );
  OR2X1 U2427 ( .IN1(n10120), .IN2(n10121), .Q(n10119) );
  AO221X1 U2428 ( .IN1(\U495/DATA1_7 ), .IN2(n14378), .IN3(\U500/DATA1_7 ), 
        .IN4(n14368), .IN5(n10122), .Q(n10121) );
  AO22X1 U2429 ( .IN1(\U470/DATA1_7 ), .IN2(n14256), .IN3(\U500/DATA2_7 ), 
        .IN4(n14356), .Q(n10122) );
  AO221X1 U2430 ( .IN1(\U475/DATA1_7 ), .IN2(n14347), .IN3(\U490/DATA1_7 ), 
        .IN4(n14335), .IN5(n10123), .Q(n10120) );
  AO22X1 U2431 ( .IN1(\U480/DATA1_7 ), .IN2(n14331), .IN3(\U485/DATA1_7 ), 
        .IN4(n14315), .Q(n10123) );
  AO221X1 U2432 ( .IN1(n5804), .IN2(n14235), .IN3(\U455/DATA1_6 ), .IN4(n14198), .IN5(n10124), .Q(n13334) );
  AO222X1 U2433 ( .IN1(\U460/DATA1_6 ), .IN2(n14412), .IN3(n14405), .IN4(
        n10125), .IN5(\U465/DATA1_6 ), .IN6(n14392), .Q(n10124) );
  OR2X1 U2434 ( .IN1(n10126), .IN2(n10127), .Q(n10125) );
  AO221X1 U2435 ( .IN1(\U495/DATA1_6 ), .IN2(n14378), .IN3(\U500/DATA1_6 ), 
        .IN4(n14369), .IN5(n10128), .Q(n10127) );
  AO22X1 U2436 ( .IN1(\U470/DATA1_6 ), .IN2(n14191), .IN3(\U500/DATA2_6 ), 
        .IN4(n14356), .Q(n10128) );
  AO221X1 U2437 ( .IN1(\U475/DATA1_6 ), .IN2(n14347), .IN3(\U490/DATA1_6 ), 
        .IN4(n14335), .IN5(n10129), .Q(n10126) );
  AO22X1 U2438 ( .IN1(\U480/DATA1_6 ), .IN2(n14326), .IN3(\U485/DATA1_6 ), 
        .IN4(n14315), .Q(n10129) );
  AO221X1 U2439 ( .IN1(n5803), .IN2(n14239), .IN3(\U455/DATA1_5 ), .IN4(n14199), .IN5(n10130), .Q(n13335) );
  AO222X1 U2440 ( .IN1(\U460/DATA1_5 ), .IN2(n14412), .IN3(n14405), .IN4(
        n10131), .IN5(\U465/DATA1_5 ), .IN6(n14392), .Q(n10130) );
  OR2X1 U2441 ( .IN1(n10132), .IN2(n10133), .Q(n10131) );
  AO221X1 U2442 ( .IN1(\U495/DATA1_5 ), .IN2(n14378), .IN3(\U500/DATA1_5 ), 
        .IN4(n14370), .IN5(n10134), .Q(n10133) );
  AO22X1 U2443 ( .IN1(\U470/DATA1_5 ), .IN2(n14190), .IN3(\U500/DATA2_5 ), 
        .IN4(n14356), .Q(n10134) );
  AO221X1 U2444 ( .IN1(\U475/DATA1_5 ), .IN2(n14347), .IN3(\U490/DATA1_5 ), 
        .IN4(n14335), .IN5(n10135), .Q(n10132) );
  AO22X1 U2445 ( .IN1(\U480/DATA1_5 ), .IN2(n14326), .IN3(\U485/DATA1_5 ), 
        .IN4(n14315), .Q(n10135) );
  AO221X1 U2446 ( .IN1(n5802), .IN2(n14240), .IN3(\U455/DATA1_4 ), .IN4(n14199), .IN5(n10136), .Q(n13336) );
  AO222X1 U2447 ( .IN1(\U460/DATA1_4 ), .IN2(n14412), .IN3(n14405), .IN4(
        n10137), .IN5(\U465/DATA1_4 ), .IN6(n14392), .Q(n10136) );
  OR2X1 U2448 ( .IN1(n10138), .IN2(n10139), .Q(n10137) );
  AO221X1 U2449 ( .IN1(\U495/DATA1_4 ), .IN2(n14378), .IN3(\U500/DATA1_4 ), 
        .IN4(n14365), .IN5(n10140), .Q(n10139) );
  AO22X1 U2450 ( .IN1(\U470/DATA1_4 ), .IN2(n14193), .IN3(\U500/DATA2_4 ), 
        .IN4(n14356), .Q(n10140) );
  AO221X1 U2451 ( .IN1(\U475/DATA1_4 ), .IN2(n14347), .IN3(\U490/DATA1_4 ), 
        .IN4(n14335), .IN5(n10141), .Q(n10138) );
  AO22X1 U2452 ( .IN1(\U480/DATA1_4 ), .IN2(n14328), .IN3(\U485/DATA1_4 ), 
        .IN4(n14315), .Q(n10141) );
  AO221X1 U2453 ( .IN1(n5801), .IN2(n14240), .IN3(\U455/DATA1_3 ), .IN4(n14199), .IN5(n10142), .Q(n13337) );
  AO222X1 U2454 ( .IN1(\U460/DATA1_3 ), .IN2(n14412), .IN3(n14405), .IN4(
        n10143), .IN5(\U465/DATA1_3 ), .IN6(n14392), .Q(n10142) );
  OR2X1 U2455 ( .IN1(n10144), .IN2(n10145), .Q(n10143) );
  AO221X1 U2456 ( .IN1(\U495/DATA1_3 ), .IN2(n14378), .IN3(\U500/DATA1_3 ), 
        .IN4(n14365), .IN5(n10146), .Q(n10145) );
  AO22X1 U2457 ( .IN1(\U470/DATA1_3 ), .IN2(n14186), .IN3(\U500/DATA2_3 ), 
        .IN4(n14356), .Q(n10146) );
  AO221X1 U2458 ( .IN1(\U475/DATA1_3 ), .IN2(n14347), .IN3(\U490/DATA1_3 ), 
        .IN4(n14335), .IN5(n10147), .Q(n10144) );
  AO22X1 U2459 ( .IN1(\U480/DATA1_3 ), .IN2(n14324), .IN3(\U485/DATA1_3 ), 
        .IN4(n14315), .Q(n10147) );
  AO221X1 U2460 ( .IN1(n5800), .IN2(n14249), .IN3(\U455/DATA1_2 ), .IN4(n14199), .IN5(n10148), .Q(n13338) );
  AO222X1 U2461 ( .IN1(\U460/DATA1_2 ), .IN2(n14413), .IN3(n14405), .IN4(
        n10149), .IN5(\U465/DATA1_2 ), .IN6(n14392), .Q(n10148) );
  OR2X1 U2462 ( .IN1(n10150), .IN2(n10151), .Q(n10149) );
  AO221X1 U2463 ( .IN1(\U495/DATA1_2 ), .IN2(n14378), .IN3(\U500/DATA1_2 ), 
        .IN4(n14364), .IN5(n10152), .Q(n10151) );
  AO22X1 U2464 ( .IN1(\U470/DATA1_2 ), .IN2(n14254), .IN3(\U500/DATA2_2 ), 
        .IN4(n14356), .Q(n10152) );
  AO221X1 U2465 ( .IN1(\U475/DATA1_2 ), .IN2(n14347), .IN3(\U490/DATA1_2 ), 
        .IN4(n14335), .IN5(n10153), .Q(n10150) );
  AO22X1 U2466 ( .IN1(\U480/DATA1_2 ), .IN2(n14326), .IN3(\U485/DATA1_2 ), 
        .IN4(n14315), .Q(n10153) );
  AO221X1 U2467 ( .IN1(n5799), .IN2(n14238), .IN3(\U455/DATA1_1 ), .IN4(n14199), .IN5(n10154), .Q(n13339) );
  AO222X1 U2468 ( .IN1(\U460/DATA1_1 ), .IN2(n14413), .IN3(n14405), .IN4(
        n10155), .IN5(\U465/DATA1_1 ), .IN6(n14392), .Q(n10154) );
  OR2X1 U2469 ( .IN1(n10156), .IN2(n10157), .Q(n10155) );
  AO221X1 U2470 ( .IN1(\U495/DATA1_1 ), .IN2(n14378), .IN3(\U500/DATA1_1 ), 
        .IN4(n14372), .IN5(n10158), .Q(n10157) );
  AO22X1 U2471 ( .IN1(\U470/DATA1_1 ), .IN2(n14257), .IN3(\U500/DATA2_1 ), 
        .IN4(n14356), .Q(n10158) );
  AO221X1 U2472 ( .IN1(\U475/DATA1_1 ), .IN2(n14347), .IN3(\U490/DATA1_1 ), 
        .IN4(n14335), .IN5(n10159), .Q(n10156) );
  AO22X1 U2473 ( .IN1(\U480/DATA1_1 ), .IN2(n14327), .IN3(\U485/DATA1_1 ), 
        .IN4(n14315), .Q(n10159) );
  AO221X1 U2474 ( .IN1(n5798), .IN2(n14239), .IN3(\U455/DATA1_0 ), .IN4(n14199), .IN5(n10160), .Q(n13340) );
  AO222X1 U2475 ( .IN1(\U460/DATA1_0 ), .IN2(n14413), .IN3(n14405), .IN4(
        n10161), .IN5(\U465/DATA1_0 ), .IN6(n14392), .Q(n10160) );
  OR2X1 U2476 ( .IN1(n10162), .IN2(n10163), .Q(n10161) );
  AO221X1 U2477 ( .IN1(\U495/DATA1_0 ), .IN2(n14378), .IN3(\U500/DATA1_0 ), 
        .IN4(n14374), .IN5(n10164), .Q(n10163) );
  AO22X1 U2478 ( .IN1(\U470/DATA1_0 ), .IN2(n14186), .IN3(\U500/DATA2_0 ), 
        .IN4(n14356), .Q(n10164) );
  AO221X1 U2479 ( .IN1(\U475/DATA1_0 ), .IN2(n14347), .IN3(\U490/DATA1_0 ), 
        .IN4(n14335), .IN5(n10165), .Q(n10162) );
  AO22X1 U2480 ( .IN1(\U480/DATA1_0 ), .IN2(n14329), .IN3(\U485/DATA1_0 ), 
        .IN4(n14315), .Q(n10165) );
  AO21X1 U2481 ( .IN1(n14240), .IN2(n13757), .IN3(n9529), .Q(n13341) );
  AO21X1 U2482 ( .IN1(n14240), .IN2(n13610), .IN3(n9531), .Q(n13342) );
  AO21X1 U2483 ( .IN1(n14240), .IN2(n14069), .IN3(n9533), .Q(n13343) );
  AO21X1 U2485 ( .IN1(n5818), .IN2(n14245), .IN3(n9534), .Q(n13344) );
  AO21X1 U2486 ( .IN1(n5817), .IN2(n14244), .IN3(n9535), .Q(n13345) );
  AO21X1 U2487 ( .IN1(n5816), .IN2(n14250), .IN3(n9536), .Q(n13346) );
  AO21X1 U2488 ( .IN1(n5815), .IN2(n14235), .IN3(n9537), .Q(n13347) );
  AO21X1 U2489 ( .IN1(n5814), .IN2(n14905), .IN3(n9538), .Q(n13348) );
  AO21X1 U2490 ( .IN1(n5813), .IN2(n14245), .IN3(n9540), .Q(n13349) );
  AO21X1 U2491 ( .IN1(n5812), .IN2(n14245), .IN3(n9542), .Q(n13350) );
  AO21X1 U2492 ( .IN1(n5811), .IN2(n14245), .IN3(n9544), .Q(n13351) );
  AO221X1 U2494 ( .IN1(n14237), .IN2(n13909), .IN3(\U508/DATA1_11 ), .IN4(
        n14199), .IN5(n10170), .Q(n13353) );
  AO222X1 U2495 ( .IN1(\U513/DATA1_11 ), .IN2(n14413), .IN3(n14395), .IN4(
        n10171), .IN5(\U518/DATA1_11 ), .IN6(n14393), .Q(n10170) );
  OR2X1 U2496 ( .IN1(n10172), .IN2(n10173), .Q(n10171) );
  AO221X1 U2497 ( .IN1(\U548/DATA1_11 ), .IN2(n14377), .IN3(\U553/DATA1_11 ), 
        .IN4(n14365), .IN5(n10174), .Q(n10173) );
  AO22X1 U2498 ( .IN1(\U523/DATA1_11 ), .IN2(n14914), .IN3(\U553/DATA2_11 ), 
        .IN4(n14356), .Q(n10174) );
  AO221X1 U2499 ( .IN1(\U528/DATA1_11 ), .IN2(n14346), .IN3(\U543/DATA1_11 ), 
        .IN4(n14334), .IN5(n10175), .Q(n10172) );
  AO22X1 U2500 ( .IN1(\U533/DATA1_11 ), .IN2(n14326), .IN3(\U538/DATA1_11 ), 
        .IN4(n14314), .Q(n10175) );
  AO221X1 U2502 ( .IN1(n14237), .IN2(n13899), .IN3(\U508/DATA1_10 ), .IN4(
        n14199), .IN5(n10177), .Q(n13354) );
  AO222X1 U2503 ( .IN1(\U513/DATA1_10 ), .IN2(n14413), .IN3(n14396), .IN4(
        n10178), .IN5(\U518/DATA1_10 ), .IN6(n14394), .Q(n10177) );
  OR2X1 U2504 ( .IN1(n10179), .IN2(n10180), .Q(n10178) );
  AO221X1 U2505 ( .IN1(\U548/DATA1_10 ), .IN2(n14377), .IN3(\U553/DATA1_10 ), 
        .IN4(n14365), .IN5(n10181), .Q(n10180) );
  AO22X1 U2506 ( .IN1(\U523/DATA1_10 ), .IN2(n14186), .IN3(\U553/DATA2_10 ), 
        .IN4(n14356), .Q(n10181) );
  AO221X1 U2507 ( .IN1(\U528/DATA1_10 ), .IN2(n14346), .IN3(\U543/DATA1_10 ), 
        .IN4(n14334), .IN5(n10182), .Q(n10179) );
  AO22X1 U2508 ( .IN1(\U533/DATA1_10 ), .IN2(n14326), .IN3(\U538/DATA1_10 ), 
        .IN4(n14314), .Q(n10182) );
  AO221X1 U2509 ( .IN1(n14236), .IN2(n14041), .IN3(\U508/DATA1_9 ), .IN4(
        n14199), .IN5(n10184), .Q(n13355) );
  AO222X1 U2510 ( .IN1(\U513/DATA1_9 ), .IN2(n14413), .IN3(n9441), .IN4(n10185), .IN5(\U518/DATA1_9 ), .IN6(n14394), .Q(n10184) );
  OR2X1 U2511 ( .IN1(n10186), .IN2(n10187), .Q(n10185) );
  AO221X1 U2512 ( .IN1(\U548/DATA1_9 ), .IN2(n14377), .IN3(\U553/DATA1_9 ), 
        .IN4(n14365), .IN5(n10188), .Q(n10187) );
  AO22X1 U2513 ( .IN1(\U523/DATA1_9 ), .IN2(n14914), .IN3(\U553/DATA2_9 ), 
        .IN4(n14356), .Q(n10188) );
  AO221X1 U2514 ( .IN1(\U528/DATA1_9 ), .IN2(n14346), .IN3(\U543/DATA1_9 ), 
        .IN4(n14334), .IN5(n10189), .Q(n10186) );
  AO22X1 U2515 ( .IN1(\U533/DATA1_9 ), .IN2(n14326), .IN3(\U538/DATA1_9 ), 
        .IN4(n14314), .Q(n10189) );
  AO221X1 U2517 ( .IN1(n5878), .IN2(n14248), .IN3(\U508/DATA1_8 ), .IN4(n14199), .IN5(n10190), .Q(n13356) );
  AO222X1 U2518 ( .IN1(\U513/DATA1_8 ), .IN2(n14413), .IN3(n14400), .IN4(
        n10191), .IN5(\U518/DATA1_8 ), .IN6(n9443), .Q(n10190) );
  OR2X1 U2519 ( .IN1(n10192), .IN2(n10193), .Q(n10191) );
  AO221X1 U2520 ( .IN1(\U548/DATA1_8 ), .IN2(n14377), .IN3(\U553/DATA1_8 ), 
        .IN4(n14365), .IN5(n10194), .Q(n10193) );
  AO22X1 U2521 ( .IN1(\U523/DATA1_8 ), .IN2(n14191), .IN3(\U553/DATA2_8 ), 
        .IN4(n14356), .Q(n10194) );
  AO221X1 U2522 ( .IN1(\U528/DATA1_8 ), .IN2(n14346), .IN3(\U543/DATA1_8 ), 
        .IN4(n14334), .IN5(n10195), .Q(n10192) );
  AO22X1 U2523 ( .IN1(\U533/DATA1_8 ), .IN2(n14326), .IN3(\U538/DATA1_8 ), 
        .IN4(n14314), .Q(n10195) );
  AO221X1 U2524 ( .IN1(n5877), .IN2(n14248), .IN3(\U508/DATA1_7 ), .IN4(n14199), .IN5(n10196), .Q(n13357) );
  AO222X1 U2525 ( .IN1(\U513/DATA1_7 ), .IN2(n14413), .IN3(n14401), .IN4(
        n10197), .IN5(\U518/DATA1_7 ), .IN6(n9443), .Q(n10196) );
  OR2X1 U2526 ( .IN1(n10198), .IN2(n10199), .Q(n10197) );
  AO221X1 U2527 ( .IN1(\U548/DATA1_7 ), .IN2(n14377), .IN3(\U553/DATA1_7 ), 
        .IN4(n14365), .IN5(n10200), .Q(n10199) );
  AO22X1 U2528 ( .IN1(\U523/DATA1_7 ), .IN2(n14254), .IN3(\U553/DATA2_7 ), 
        .IN4(n14356), .Q(n10200) );
  AO221X1 U2529 ( .IN1(\U528/DATA1_7 ), .IN2(n14346), .IN3(\U543/DATA1_7 ), 
        .IN4(n14334), .IN5(n10201), .Q(n10198) );
  AO22X1 U2530 ( .IN1(\U533/DATA1_7 ), .IN2(n14326), .IN3(\U538/DATA1_7 ), 
        .IN4(n14314), .Q(n10201) );
  AO221X1 U2531 ( .IN1(n5876), .IN2(n14248), .IN3(\U508/DATA1_6 ), .IN4(n14199), .IN5(n10202), .Q(n13358) );
  AO222X1 U2532 ( .IN1(\U513/DATA1_6 ), .IN2(n14413), .IN3(n14402), .IN4(
        n10203), .IN5(\U518/DATA1_6 ), .IN6(n9443), .Q(n10202) );
  OR2X1 U2533 ( .IN1(n10204), .IN2(n10205), .Q(n10203) );
  AO221X1 U2534 ( .IN1(\U548/DATA1_6 ), .IN2(n14377), .IN3(\U553/DATA1_6 ), 
        .IN4(n14365), .IN5(n10206), .Q(n10205) );
  AO22X1 U2535 ( .IN1(\U523/DATA1_6 ), .IN2(n14257), .IN3(\U553/DATA2_6 ), 
        .IN4(n14356), .Q(n10206) );
  AO221X1 U2536 ( .IN1(\U528/DATA1_6 ), .IN2(n14346), .IN3(\U543/DATA1_6 ), 
        .IN4(n14334), .IN5(n10207), .Q(n10204) );
  AO22X1 U2537 ( .IN1(\U533/DATA1_6 ), .IN2(n14326), .IN3(\U538/DATA1_6 ), 
        .IN4(n14314), .Q(n10207) );
  AO221X1 U2538 ( .IN1(n5875), .IN2(n14248), .IN3(\U508/DATA1_5 ), .IN4(n14200), .IN5(n10208), .Q(n13359) );
  AO222X1 U2539 ( .IN1(\U513/DATA1_5 ), .IN2(n14413), .IN3(n14403), .IN4(
        n10209), .IN5(\U518/DATA1_5 ), .IN6(n9443), .Q(n10208) );
  OR2X1 U2540 ( .IN1(n10210), .IN2(n10211), .Q(n10209) );
  AO221X1 U2541 ( .IN1(\U548/DATA1_5 ), .IN2(n14377), .IN3(\U553/DATA1_5 ), 
        .IN4(n14365), .IN5(n10212), .Q(n10211) );
  AO22X1 U2542 ( .IN1(\U523/DATA1_5 ), .IN2(n14255), .IN3(\U553/DATA2_5 ), 
        .IN4(n14356), .Q(n10212) );
  AO221X1 U2543 ( .IN1(\U528/DATA1_5 ), .IN2(n14346), .IN3(\U543/DATA1_5 ), 
        .IN4(n14334), .IN5(n10213), .Q(n10210) );
  AO22X1 U2544 ( .IN1(\U533/DATA1_5 ), .IN2(n14326), .IN3(\U538/DATA1_5 ), 
        .IN4(n14314), .Q(n10213) );
  AO221X1 U2545 ( .IN1(n5874), .IN2(n14248), .IN3(\U508/DATA1_4 ), .IN4(n14200), .IN5(n10214), .Q(n13360) );
  AO222X1 U2546 ( .IN1(\U513/DATA1_4 ), .IN2(n14413), .IN3(n14402), .IN4(
        n10215), .IN5(\U518/DATA1_4 ), .IN6(n14390), .Q(n10214) );
  OR2X1 U2547 ( .IN1(n10216), .IN2(n10217), .Q(n10215) );
  AO221X1 U2548 ( .IN1(\U548/DATA1_4 ), .IN2(n14377), .IN3(\U553/DATA1_4 ), 
        .IN4(n14365), .IN5(n10218), .Q(n10217) );
  AO22X1 U2549 ( .IN1(\U523/DATA1_4 ), .IN2(n14255), .IN3(\U553/DATA2_4 ), 
        .IN4(n14355), .Q(n10218) );
  AO221X1 U2550 ( .IN1(\U528/DATA1_4 ), .IN2(n14346), .IN3(\U543/DATA1_4 ), 
        .IN4(n14334), .IN5(n10219), .Q(n10216) );
  AO22X1 U2551 ( .IN1(\U533/DATA1_4 ), .IN2(n14326), .IN3(\U538/DATA1_4 ), 
        .IN4(n14314), .Q(n10219) );
  AO221X1 U2552 ( .IN1(n5873), .IN2(n14248), .IN3(\U508/DATA1_3 ), .IN4(n14200), .IN5(n10220), .Q(n13361) );
  AO222X1 U2553 ( .IN1(\U513/DATA1_3 ), .IN2(n14413), .IN3(n14404), .IN4(
        n10221), .IN5(\U518/DATA1_3 ), .IN6(n9443), .Q(n10220) );
  OR2X1 U2554 ( .IN1(n10222), .IN2(n10223), .Q(n10221) );
  AO221X1 U2555 ( .IN1(\U548/DATA1_3 ), .IN2(n14377), .IN3(\U553/DATA1_3 ), 
        .IN4(n14365), .IN5(n10224), .Q(n10223) );
  AO22X1 U2556 ( .IN1(\U523/DATA1_3 ), .IN2(n14191), .IN3(\U553/DATA2_3 ), 
        .IN4(n14355), .Q(n10224) );
  AO221X1 U2557 ( .IN1(\U528/DATA1_3 ), .IN2(n14346), .IN3(\U543/DATA1_3 ), 
        .IN4(n14334), .IN5(n10225), .Q(n10222) );
  AO22X1 U2558 ( .IN1(\U533/DATA1_3 ), .IN2(n14326), .IN3(\U538/DATA1_3 ), 
        .IN4(n14314), .Q(n10225) );
  AO221X1 U2559 ( .IN1(n5872), .IN2(n14247), .IN3(\U508/DATA1_2 ), .IN4(n14200), .IN5(n10226), .Q(n13362) );
  AO222X1 U2560 ( .IN1(\U513/DATA1_2 ), .IN2(n14413), .IN3(n14405), .IN4(
        n10227), .IN5(\U518/DATA1_2 ), .IN6(n14389), .Q(n10226) );
  OR2X1 U2561 ( .IN1(n10228), .IN2(n10229), .Q(n10227) );
  AO221X1 U2562 ( .IN1(\U548/DATA1_2 ), .IN2(n14377), .IN3(\U553/DATA1_2 ), 
        .IN4(n14365), .IN5(n10230), .Q(n10229) );
  AO22X1 U2563 ( .IN1(\U523/DATA1_2 ), .IN2(n14256), .IN3(\U553/DATA2_2 ), 
        .IN4(n14355), .Q(n10230) );
  AO221X1 U2564 ( .IN1(\U528/DATA1_2 ), .IN2(n14346), .IN3(\U543/DATA1_2 ), 
        .IN4(n14334), .IN5(n10231), .Q(n10228) );
  AO22X1 U2565 ( .IN1(\U533/DATA1_2 ), .IN2(n14326), .IN3(\U538/DATA1_2 ), 
        .IN4(n14314), .Q(n10231) );
  AO221X1 U2566 ( .IN1(n5871), .IN2(n14247), .IN3(\U508/DATA1_1 ), .IN4(n14200), .IN5(n10232), .Q(n13363) );
  AO222X1 U2567 ( .IN1(\U513/DATA1_1 ), .IN2(n14413), .IN3(n14396), .IN4(
        n10233), .IN5(\U518/DATA1_1 ), .IN6(n14390), .Q(n10232) );
  OR2X1 U2568 ( .IN1(n10234), .IN2(n10235), .Q(n10233) );
  AO221X1 U2569 ( .IN1(\U548/DATA1_1 ), .IN2(n14377), .IN3(\U553/DATA1_1 ), 
        .IN4(n14365), .IN5(n10236), .Q(n10235) );
  AO22X1 U2570 ( .IN1(\U523/DATA1_1 ), .IN2(n14186), .IN3(\U553/DATA2_1 ), 
        .IN4(n14355), .Q(n10236) );
  AO221X1 U2571 ( .IN1(\U528/DATA1_1 ), .IN2(n14346), .IN3(\U543/DATA1_1 ), 
        .IN4(n14334), .IN5(n10237), .Q(n10234) );
  AO22X1 U2572 ( .IN1(\U533/DATA1_1 ), .IN2(n14326), .IN3(\U538/DATA1_1 ), 
        .IN4(n14314), .Q(n10237) );
  AO221X1 U2573 ( .IN1(n5870), .IN2(n14247), .IN3(\U508/DATA1_0 ), .IN4(n14200), .IN5(n10238), .Q(n13364) );
  AO222X1 U2574 ( .IN1(\U513/DATA1_0 ), .IN2(n14413), .IN3(n9441), .IN4(n10239), .IN5(\U518/DATA1_0 ), .IN6(n14391), .Q(n10238) );
  OR2X1 U2575 ( .IN1(n10240), .IN2(n10241), .Q(n10239) );
  AO221X1 U2576 ( .IN1(\U548/DATA1_0 ), .IN2(n14377), .IN3(\U553/DATA1_0 ), 
        .IN4(n14365), .IN5(n10242), .Q(n10241) );
  AO22X1 U2577 ( .IN1(\U523/DATA1_0 ), .IN2(n14254), .IN3(\U553/DATA2_0 ), 
        .IN4(n14355), .Q(n10242) );
  AO221X1 U2578 ( .IN1(\U528/DATA1_0 ), .IN2(n14346), .IN3(\U543/DATA1_0 ), 
        .IN4(n14334), .IN5(n10243), .Q(n10240) );
  AO22X1 U2579 ( .IN1(\U533/DATA1_0 ), .IN2(n14326), .IN3(\U538/DATA1_0 ), 
        .IN4(n14314), .Q(n10243) );
  AO21X1 U2580 ( .IN1(n14239), .IN2(n13756), .IN3(n9529), .Q(n13365) );
  AO21X1 U2581 ( .IN1(n14239), .IN2(n13609), .IN3(n9531), .Q(n13366) );
  AO21X1 U2582 ( .IN1(n14239), .IN2(n14068), .IN3(n9533), .Q(n13367) );
  AO21X1 U2584 ( .IN1(n5890), .IN2(n14245), .IN3(n9534), .Q(n13368) );
  AO21X1 U2585 ( .IN1(n5889), .IN2(n14245), .IN3(n9535), .Q(n13369) );
  AO21X1 U2586 ( .IN1(n5888), .IN2(n14245), .IN3(n9536), .Q(n13370) );
  AO21X1 U2587 ( .IN1(n5887), .IN2(n14245), .IN3(n9537), .Q(n13371) );
  AO21X1 U2588 ( .IN1(n5886), .IN2(n14245), .IN3(n9538), .Q(n13372) );
  AO21X1 U2589 ( .IN1(n5885), .IN2(n14245), .IN3(n9540), .Q(n13373) );
  AO21X1 U2590 ( .IN1(n5884), .IN2(n14245), .IN3(n9542), .Q(n13374) );
  AO21X1 U2591 ( .IN1(n5883), .IN2(n14245), .IN3(n9544), .Q(n13375) );
  AO221X1 U2592 ( .IN1(n14236), .IN2(n13908), .IN3(\U570/DATA1_11 ), .IN4(
        n14200), .IN5(n10248), .Q(n13376) );
  AO222X1 U2593 ( .IN1(\U575/DATA1_11 ), .IN2(n14414), .IN3(n14397), .IN4(
        n10249), .IN5(\U580/DATA1_11 ), .IN6(n14393), .Q(n10248) );
  OR2X1 U2594 ( .IN1(n10250), .IN2(n10251), .Q(n10249) );
  AO221X1 U2595 ( .IN1(\U610/DATA1_11 ), .IN2(n14376), .IN3(\U615/DATA1_11 ), 
        .IN4(n14364), .IN5(n10252), .Q(n10251) );
  AO22X1 U2596 ( .IN1(\U585/DATA1_11 ), .IN2(n14191), .IN3(\U615/DATA2_11 ), 
        .IN4(n14355), .Q(n10252) );
  AO221X1 U2597 ( .IN1(\U590/DATA1_11 ), .IN2(n14345), .IN3(\U605/DATA1_11 ), 
        .IN4(n14334), .IN5(n10253), .Q(n10250) );
  AO22X1 U2598 ( .IN1(\U595/DATA1_11 ), .IN2(n14325), .IN3(\U600/DATA1_11 ), 
        .IN4(n14313), .Q(n10253) );
  AO221X1 U2600 ( .IN1(n14236), .IN2(n13898), .IN3(\U570/DATA1_10 ), .IN4(
        n14258), .IN5(n10255), .Q(n13377) );
  AO222X1 U2601 ( .IN1(\U575/DATA1_10 ), .IN2(n14414), .IN3(n14398), .IN4(
        n10256), .IN5(\U580/DATA1_10 ), .IN6(n14393), .Q(n10255) );
  OR2X1 U2602 ( .IN1(n10257), .IN2(n10258), .Q(n10256) );
  AO221X1 U2603 ( .IN1(\U610/DATA1_10 ), .IN2(n14376), .IN3(\U615/DATA1_10 ), 
        .IN4(n14364), .IN5(n10259), .Q(n10258) );
  AO22X1 U2604 ( .IN1(\U585/DATA1_10 ), .IN2(n14192), .IN3(\U615/DATA2_10 ), 
        .IN4(n14355), .Q(n10259) );
  AO221X1 U2605 ( .IN1(\U590/DATA1_10 ), .IN2(n14345), .IN3(\U605/DATA1_10 ), 
        .IN4(n14340), .IN5(n10260), .Q(n10257) );
  AO22X1 U2606 ( .IN1(\U595/DATA1_10 ), .IN2(n14325), .IN3(\U600/DATA1_10 ), 
        .IN4(n14313), .Q(n10260) );
  AO221X1 U2607 ( .IN1(n14236), .IN2(n14040), .IN3(\U570/DATA1_9 ), .IN4(
        n14258), .IN5(n10262), .Q(n13378) );
  AO222X1 U2608 ( .IN1(\U575/DATA1_9 ), .IN2(n14414), .IN3(n14399), .IN4(
        n10263), .IN5(\U580/DATA1_9 ), .IN6(n14393), .Q(n10262) );
  OR2X1 U2609 ( .IN1(n10264), .IN2(n10265), .Q(n10263) );
  AO221X1 U2610 ( .IN1(\U610/DATA1_9 ), .IN2(n14376), .IN3(\U615/DATA1_9 ), 
        .IN4(n14364), .IN5(n10266), .Q(n10265) );
  AO22X1 U2611 ( .IN1(\U585/DATA1_9 ), .IN2(n14256), .IN3(\U615/DATA2_9 ), 
        .IN4(n14355), .Q(n10266) );
  AO221X1 U2612 ( .IN1(\U590/DATA1_9 ), .IN2(n14345), .IN3(\U605/DATA1_9 ), 
        .IN4(n14343), .IN5(n10267), .Q(n10264) );
  AO22X1 U2613 ( .IN1(\U595/DATA1_9 ), .IN2(n14325), .IN3(\U600/DATA1_9 ), 
        .IN4(n14313), .Q(n10267) );
  AO221X1 U2615 ( .IN1(n5950), .IN2(n14249), .IN3(\U570/DATA1_8 ), .IN4(n14258), .IN5(n10268), .Q(n13379) );
  AO222X1 U2616 ( .IN1(\U575/DATA1_8 ), .IN2(n14414), .IN3(n14395), .IN4(
        n10269), .IN5(\U580/DATA1_8 ), .IN6(n14393), .Q(n10268) );
  OR2X1 U2617 ( .IN1(n10270), .IN2(n10271), .Q(n10269) );
  AO221X1 U2618 ( .IN1(\U610/DATA1_8 ), .IN2(n14376), .IN3(\U615/DATA1_8 ), 
        .IN4(n14364), .IN5(n10272), .Q(n10271) );
  AO22X1 U2619 ( .IN1(\U585/DATA1_8 ), .IN2(n14189), .IN3(\U615/DATA2_8 ), 
        .IN4(n14355), .Q(n10272) );
  AO221X1 U2620 ( .IN1(\U590/DATA1_8 ), .IN2(n14345), .IN3(\U605/DATA1_8 ), 
        .IN4(n14336), .IN5(n10273), .Q(n10270) );
  AO22X1 U2621 ( .IN1(\U595/DATA1_8 ), .IN2(n14325), .IN3(\U600/DATA1_8 ), 
        .IN4(n14313), .Q(n10273) );
  AO221X1 U2622 ( .IN1(n5949), .IN2(n14248), .IN3(\U570/DATA1_7 ), .IN4(n14258), .IN5(n10274), .Q(n13380) );
  AO222X1 U2623 ( .IN1(\U575/DATA1_7 ), .IN2(n14414), .IN3(n14403), .IN4(
        n10275), .IN5(\U580/DATA1_7 ), .IN6(n14393), .Q(n10274) );
  OR2X1 U2624 ( .IN1(n10276), .IN2(n10277), .Q(n10275) );
  AO221X1 U2625 ( .IN1(\U610/DATA1_7 ), .IN2(n14376), .IN3(\U615/DATA1_7 ), 
        .IN4(n14364), .IN5(n10278), .Q(n10277) );
  AO22X1 U2626 ( .IN1(\U585/DATA1_7 ), .IN2(n14193), .IN3(\U615/DATA2_7 ), 
        .IN4(n14355), .Q(n10278) );
  AO221X1 U2627 ( .IN1(\U590/DATA1_7 ), .IN2(n14345), .IN3(\U605/DATA1_7 ), 
        .IN4(n14337), .IN5(n10279), .Q(n10276) );
  AO22X1 U2628 ( .IN1(\U595/DATA1_7 ), .IN2(n14325), .IN3(\U600/DATA1_7 ), 
        .IN4(n14313), .Q(n10279) );
  AO221X1 U2629 ( .IN1(n5948), .IN2(n14247), .IN3(\U570/DATA1_6 ), .IN4(n14258), .IN5(n10280), .Q(n13381) );
  AO222X1 U2630 ( .IN1(\U575/DATA1_6 ), .IN2(n14414), .IN3(n14404), .IN4(
        n10281), .IN5(\U580/DATA1_6 ), .IN6(n14393), .Q(n10280) );
  OR2X1 U2631 ( .IN1(n10282), .IN2(n10283), .Q(n10281) );
  AO221X1 U2632 ( .IN1(\U610/DATA1_6 ), .IN2(n14376), .IN3(\U615/DATA1_6 ), 
        .IN4(n14364), .IN5(n10284), .Q(n10283) );
  AO22X1 U2633 ( .IN1(\U585/DATA1_6 ), .IN2(n14914), .IN3(\U615/DATA2_6 ), 
        .IN4(n14355), .Q(n10284) );
  AO221X1 U2634 ( .IN1(\U590/DATA1_6 ), .IN2(n14345), .IN3(\U605/DATA1_6 ), 
        .IN4(n14338), .IN5(n10285), .Q(n10282) );
  AO22X1 U2635 ( .IN1(\U595/DATA1_6 ), .IN2(n14325), .IN3(\U600/DATA1_6 ), 
        .IN4(n14313), .Q(n10285) );
  AO221X1 U2636 ( .IN1(n5947), .IN2(n14242), .IN3(\U570/DATA1_5 ), .IN4(n14258), .IN5(n10286), .Q(n13382) );
  AO222X1 U2637 ( .IN1(\U575/DATA1_5 ), .IN2(n14414), .IN3(n14405), .IN4(
        n10287), .IN5(\U580/DATA1_5 ), .IN6(n14393), .Q(n10286) );
  OR2X1 U2638 ( .IN1(n10288), .IN2(n10289), .Q(n10287) );
  AO221X1 U2639 ( .IN1(\U610/DATA1_5 ), .IN2(n14376), .IN3(\U615/DATA1_5 ), 
        .IN4(n14364), .IN5(n10290), .Q(n10289) );
  AO22X1 U2640 ( .IN1(\U585/DATA1_5 ), .IN2(n14191), .IN3(\U615/DATA2_5 ), 
        .IN4(n14355), .Q(n10290) );
  AO221X1 U2641 ( .IN1(\U590/DATA1_5 ), .IN2(n14345), .IN3(\U605/DATA1_5 ), 
        .IN4(n14339), .IN5(n10291), .Q(n10288) );
  AO22X1 U2642 ( .IN1(\U595/DATA1_5 ), .IN2(n14325), .IN3(\U600/DATA1_5 ), 
        .IN4(n14313), .Q(n10291) );
  AO221X1 U2643 ( .IN1(n5946), .IN2(n14236), .IN3(\U570/DATA1_4 ), .IN4(n14258), .IN5(n10292), .Q(n13383) );
  AO222X1 U2644 ( .IN1(\U575/DATA1_4 ), .IN2(n14414), .IN3(n9441), .IN4(n10293), .IN5(\U580/DATA1_4 ), .IN6(n14393), .Q(n10292) );
  OR2X1 U2645 ( .IN1(n10294), .IN2(n10295), .Q(n10293) );
  AO221X1 U2646 ( .IN1(\U610/DATA1_4 ), .IN2(n14376), .IN3(\U615/DATA1_4 ), 
        .IN4(n14364), .IN5(n10296), .Q(n10295) );
  AO22X1 U2647 ( .IN1(\U585/DATA1_4 ), .IN2(n14192), .IN3(\U615/DATA2_4 ), 
        .IN4(n14355), .Q(n10296) );
  AO221X1 U2648 ( .IN1(\U590/DATA1_4 ), .IN2(n14345), .IN3(\U605/DATA1_4 ), 
        .IN4(n14334), .IN5(n10297), .Q(n10294) );
  AO22X1 U2649 ( .IN1(\U595/DATA1_4 ), .IN2(n14325), .IN3(\U600/DATA1_4 ), 
        .IN4(n14313), .Q(n10297) );
  AO221X1 U2650 ( .IN1(n5945), .IN2(n14242), .IN3(\U570/DATA1_3 ), .IN4(n14258), .IN5(n10298), .Q(n13384) );
  AO222X1 U2651 ( .IN1(\U575/DATA1_3 ), .IN2(n14414), .IN3(n14400), .IN4(
        n10299), .IN5(\U580/DATA1_3 ), .IN6(n14393), .Q(n10298) );
  OR2X1 U2652 ( .IN1(n10300), .IN2(n10301), .Q(n10299) );
  AO221X1 U2653 ( .IN1(\U610/DATA1_3 ), .IN2(n14376), .IN3(\U615/DATA1_3 ), 
        .IN4(n14364), .IN5(n10302), .Q(n10301) );
  AO22X1 U2654 ( .IN1(\U585/DATA1_3 ), .IN2(n14256), .IN3(\U615/DATA2_3 ), 
        .IN4(n14355), .Q(n10302) );
  AO221X1 U2655 ( .IN1(\U590/DATA1_3 ), .IN2(n14345), .IN3(\U605/DATA1_3 ), 
        .IN4(n14340), .IN5(n10303), .Q(n10300) );
  AO22X1 U2656 ( .IN1(\U595/DATA1_3 ), .IN2(n14325), .IN3(\U600/DATA1_3 ), 
        .IN4(n14313), .Q(n10303) );
  AO221X1 U2657 ( .IN1(n5944), .IN2(n14241), .IN3(\U570/DATA1_2 ), .IN4(n14258), .IN5(n10304), .Q(n13385) );
  AO222X1 U2658 ( .IN1(\U575/DATA1_2 ), .IN2(n14414), .IN3(n14401), .IN4(
        n10305), .IN5(\U580/DATA1_2 ), .IN6(n14393), .Q(n10304) );
  OR2X1 U2659 ( .IN1(n10306), .IN2(n10307), .Q(n10305) );
  AO221X1 U2660 ( .IN1(\U610/DATA1_2 ), .IN2(n14376), .IN3(\U615/DATA1_2 ), 
        .IN4(n14364), .IN5(n10308), .Q(n10307) );
  AO22X1 U2661 ( .IN1(\U585/DATA1_2 ), .IN2(n14254), .IN3(\U615/DATA2_2 ), 
        .IN4(n14355), .Q(n10308) );
  AO221X1 U2662 ( .IN1(\U590/DATA1_2 ), .IN2(n14345), .IN3(\U605/DATA1_2 ), 
        .IN4(n14340), .IN5(n10309), .Q(n10306) );
  AO22X1 U2663 ( .IN1(\U595/DATA1_2 ), .IN2(n14325), .IN3(\U600/DATA1_2 ), 
        .IN4(n14313), .Q(n10309) );
  AO221X1 U2664 ( .IN1(n5943), .IN2(n14241), .IN3(\U570/DATA1_1 ), .IN4(n14258), .IN5(n10310), .Q(n13386) );
  AO222X1 U2665 ( .IN1(\U575/DATA1_1 ), .IN2(n14414), .IN3(n14395), .IN4(
        n10311), .IN5(\U580/DATA1_1 ), .IN6(n14393), .Q(n10310) );
  OR2X1 U2666 ( .IN1(n10312), .IN2(n10313), .Q(n10311) );
  AO221X1 U2667 ( .IN1(\U610/DATA1_1 ), .IN2(n14376), .IN3(\U615/DATA1_1 ), 
        .IN4(n14364), .IN5(n10314), .Q(n10313) );
  AO22X1 U2668 ( .IN1(\U585/DATA1_1 ), .IN2(n14914), .IN3(\U615/DATA2_1 ), 
        .IN4(n9450), .Q(n10314) );
  AO221X1 U2669 ( .IN1(\U590/DATA1_1 ), .IN2(n14345), .IN3(\U605/DATA1_1 ), 
        .IN4(n14334), .IN5(n10315), .Q(n10312) );
  AO22X1 U2670 ( .IN1(\U595/DATA1_1 ), .IN2(n14325), .IN3(\U600/DATA1_1 ), 
        .IN4(n14313), .Q(n10315) );
  AO221X1 U2671 ( .IN1(n5942), .IN2(n14238), .IN3(\U570/DATA1_0 ), .IN4(n14258), .IN5(n10316), .Q(n13387) );
  AO222X1 U2672 ( .IN1(\U575/DATA1_0 ), .IN2(n14414), .IN3(n9441), .IN4(n10317), .IN5(\U580/DATA1_0 ), .IN6(n14393), .Q(n10316) );
  OR2X1 U2673 ( .IN1(n10318), .IN2(n10319), .Q(n10317) );
  AO221X1 U2674 ( .IN1(\U610/DATA1_0 ), .IN2(n14376), .IN3(\U615/DATA1_0 ), 
        .IN4(n14364), .IN5(n10320), .Q(n10319) );
  AO22X1 U2675 ( .IN1(\U585/DATA1_0 ), .IN2(n14254), .IN3(\U615/DATA2_0 ), 
        .IN4(n9450), .Q(n10320) );
  AO221X1 U2676 ( .IN1(\U590/DATA1_0 ), .IN2(n14345), .IN3(\U605/DATA1_0 ), 
        .IN4(n14335), .IN5(n10321), .Q(n10318) );
  AO22X1 U2677 ( .IN1(\U595/DATA1_0 ), .IN2(n14325), .IN3(\U600/DATA1_0 ), 
        .IN4(n14313), .Q(n10321) );
  AO21X1 U2678 ( .IN1(n14239), .IN2(n13755), .IN3(n9529), .Q(n13388) );
  AO22X1 U2680 ( .IN1(\U571/DATA1_11 ), .IN2(n14258), .IN3(\U581/DATA1_11 ), 
        .IN4(n14394), .Q(n10324) );
  OR2X1 U2681 ( .IN1(n10325), .IN2(n10326), .Q(n10323) );
  AO221X1 U2682 ( .IN1(\U611/DATA1_11 ), .IN2(n9446), .IN3(\U616/DATA1_11 ), 
        .IN4(n14365), .IN5(n10327), .Q(n10326) );
  AO22X1 U2683 ( .IN1(\U586/DATA1_11 ), .IN2(n14189), .IN3(\U616/DATA2_11 ), 
        .IN4(n9450), .Q(n10327) );
  AO221X1 U2684 ( .IN1(\U591/DATA1_11 ), .IN2(n9451), .IN3(\U606/DATA1_11 ), 
        .IN4(n14343), .IN5(n10328), .Q(n10325) );
  AO22X1 U2685 ( .IN1(\U596/DATA1_11 ), .IN2(n14324), .IN3(\U601/DATA1_11 ), 
        .IN4(n9455), .Q(n10328) );
  AO21X1 U2686 ( .IN1(n14238), .IN2(n13608), .IN3(n9531), .Q(n13389) );
  AO22X1 U2688 ( .IN1(\U571/DATA1_10 ), .IN2(n14258), .IN3(\U581/DATA1_10 ), 
        .IN4(n14394), .Q(n10331) );
  OR2X1 U2689 ( .IN1(n10332), .IN2(n10333), .Q(n10330) );
  AO221X1 U2690 ( .IN1(\U611/DATA1_10 ), .IN2(n9446), .IN3(\U616/DATA1_10 ), 
        .IN4(n9447), .IN5(n10334), .Q(n10333) );
  AO22X1 U2691 ( .IN1(\U586/DATA1_10 ), .IN2(n14192), .IN3(\U616/DATA2_10 ), 
        .IN4(n9450), .Q(n10334) );
  AO221X1 U2692 ( .IN1(\U591/DATA1_10 ), .IN2(n9451), .IN3(\U606/DATA1_10 ), 
        .IN4(n9452), .IN5(n10335), .Q(n10332) );
  AO22X1 U2693 ( .IN1(\U596/DATA1_10 ), .IN2(n9454), .IN3(\U601/DATA1_10 ), 
        .IN4(n9455), .Q(n10335) );
  AO21X1 U2694 ( .IN1(n14241), .IN2(n14067), .IN3(n9533), .Q(n13390) );
  AO22X1 U2696 ( .IN1(\U571/DATA1_9 ), .IN2(n14258), .IN3(\U581/DATA1_9 ), 
        .IN4(n14394), .Q(n10338) );
  OR2X1 U2697 ( .IN1(n10339), .IN2(n10340), .Q(n10337) );
  AO221X1 U2698 ( .IN1(\U611/DATA1_9 ), .IN2(n9446), .IN3(\U616/DATA1_9 ), 
        .IN4(n9447), .IN5(n10341), .Q(n10340) );
  AO22X1 U2699 ( .IN1(\U586/DATA1_9 ), .IN2(n14192), .IN3(\U616/DATA2_9 ), 
        .IN4(n9450), .Q(n10341) );
  AO221X1 U2700 ( .IN1(\U591/DATA1_9 ), .IN2(n9451), .IN3(\U606/DATA1_9 ), 
        .IN4(n9452), .IN5(n10342), .Q(n10339) );
  AO22X1 U2701 ( .IN1(\U596/DATA1_9 ), .IN2(n9454), .IN3(\U601/DATA1_9 ), 
        .IN4(n9455), .Q(n10342) );
  AO21X1 U2703 ( .IN1(n5962), .IN2(n14245), .IN3(n9534), .Q(n13391) );
  AO22X1 U2705 ( .IN1(\U571/DATA1_8 ), .IN2(n14258), .IN3(\U581/DATA1_8 ), 
        .IN4(n14394), .Q(n10344) );
  OR2X1 U2706 ( .IN1(n10345), .IN2(n10346), .Q(n10343) );
  AO221X1 U2707 ( .IN1(\U611/DATA1_8 ), .IN2(n9446), .IN3(\U616/DATA1_8 ), 
        .IN4(n14374), .IN5(n10347), .Q(n10346) );
  AO22X1 U2708 ( .IN1(\U586/DATA1_8 ), .IN2(n14257), .IN3(\U616/DATA2_8 ), 
        .IN4(n14363), .Q(n10347) );
  AO221X1 U2709 ( .IN1(\U591/DATA1_8 ), .IN2(n9451), .IN3(\U606/DATA1_8 ), 
        .IN4(n14343), .IN5(n10348), .Q(n10345) );
  AO22X1 U2710 ( .IN1(\U596/DATA1_8 ), .IN2(n9454), .IN3(\U601/DATA1_8 ), 
        .IN4(n9455), .Q(n10348) );
  AO21X1 U2711 ( .IN1(n5961), .IN2(n14245), .IN3(n9535), .Q(n13392) );
  AO22X1 U2713 ( .IN1(\U571/DATA1_7 ), .IN2(n14258), .IN3(\U581/DATA1_7 ), 
        .IN4(n14394), .Q(n10350) );
  OR2X1 U2714 ( .IN1(n10351), .IN2(n10352), .Q(n10349) );
  AO221X1 U2715 ( .IN1(\U611/DATA1_7 ), .IN2(n9446), .IN3(\U616/DATA1_7 ), 
        .IN4(n9447), .IN5(n10353), .Q(n10352) );
  AO22X1 U2716 ( .IN1(\U586/DATA1_7 ), .IN2(n14190), .IN3(\U616/DATA2_7 ), 
        .IN4(n9450), .Q(n10353) );
  AO221X1 U2717 ( .IN1(\U591/DATA1_7 ), .IN2(n9451), .IN3(\U606/DATA1_7 ), 
        .IN4(n14334), .IN5(n10354), .Q(n10351) );
  AO22X1 U2718 ( .IN1(\U596/DATA1_7 ), .IN2(n14326), .IN3(\U601/DATA1_7 ), 
        .IN4(n9455), .Q(n10354) );
  AO21X1 U2719 ( .IN1(n5960), .IN2(n14244), .IN3(n9536), .Q(n13393) );
  AO22X1 U2721 ( .IN1(\U571/DATA1_6 ), .IN2(n14258), .IN3(\U581/DATA1_6 ), 
        .IN4(n14394), .Q(n10356) );
  OR2X1 U2722 ( .IN1(n10357), .IN2(n10358), .Q(n10355) );
  AO221X1 U2723 ( .IN1(\U611/DATA1_6 ), .IN2(n9446), .IN3(\U616/DATA1_6 ), 
        .IN4(n9447), .IN5(n10359), .Q(n10358) );
  AO22X1 U2724 ( .IN1(\U586/DATA1_6 ), .IN2(n14193), .IN3(\U616/DATA2_6 ), 
        .IN4(n9450), .Q(n10359) );
  AO221X1 U2725 ( .IN1(\U591/DATA1_6 ), .IN2(n14344), .IN3(\U606/DATA1_6 ), 
        .IN4(n9452), .IN5(n10360), .Q(n10357) );
  AO22X1 U2726 ( .IN1(\U596/DATA1_6 ), .IN2(n9454), .IN3(\U601/DATA1_6 ), 
        .IN4(n9455), .Q(n10360) );
  AO21X1 U2727 ( .IN1(n5959), .IN2(n14244), .IN3(n9537), .Q(n13394) );
  AO22X1 U2729 ( .IN1(\U571/DATA1_5 ), .IN2(n14258), .IN3(\U581/DATA1_5 ), 
        .IN4(n14394), .Q(n10362) );
  OR2X1 U2730 ( .IN1(n10363), .IN2(n10364), .Q(n10361) );
  AO221X1 U2731 ( .IN1(\U611/DATA1_5 ), .IN2(n9446), .IN3(\U616/DATA1_5 ), 
        .IN4(n9447), .IN5(n10365), .Q(n10364) );
  AO22X1 U2732 ( .IN1(\U586/DATA1_5 ), .IN2(n14255), .IN3(\U616/DATA2_5 ), 
        .IN4(n9450), .Q(n10365) );
  AO221X1 U2733 ( .IN1(\U591/DATA1_5 ), .IN2(n9451), .IN3(\U606/DATA1_5 ), 
        .IN4(n14339), .IN5(n10366), .Q(n10363) );
  AO22X1 U2734 ( .IN1(\U596/DATA1_5 ), .IN2(n14324), .IN3(\U601/DATA1_5 ), 
        .IN4(n9455), .Q(n10366) );
  AO21X1 U2735 ( .IN1(n5958), .IN2(n14244), .IN3(n9538), .Q(n13395) );
  AO22X1 U2737 ( .IN1(\U571/DATA1_4 ), .IN2(n14258), .IN3(\U581/DATA1_4 ), 
        .IN4(n14394), .Q(n10368) );
  OR2X1 U2738 ( .IN1(n10369), .IN2(n10370), .Q(n10367) );
  AO221X1 U2739 ( .IN1(\U611/DATA1_4 ), .IN2(n9446), .IN3(\U616/DATA1_4 ), 
        .IN4(n9447), .IN5(n10371), .Q(n10370) );
  AO22X1 U2740 ( .IN1(\U586/DATA1_4 ), .IN2(n14190), .IN3(\U616/DATA2_4 ), 
        .IN4(n14362), .Q(n10371) );
  AO221X1 U2741 ( .IN1(\U591/DATA1_4 ), .IN2(n9451), .IN3(\U606/DATA1_4 ), 
        .IN4(n14343), .IN5(n10372), .Q(n10369) );
  AO22X1 U2742 ( .IN1(\U596/DATA1_4 ), .IN2(n9454), .IN3(\U601/DATA1_4 ), 
        .IN4(n9455), .Q(n10372) );
  AO21X1 U2743 ( .IN1(n5957), .IN2(n14244), .IN3(n9540), .Q(n13396) );
  AO22X1 U2745 ( .IN1(\U571/DATA1_3 ), .IN2(n14258), .IN3(\U581/DATA1_3 ), 
        .IN4(n14394), .Q(n10374) );
  OR2X1 U2746 ( .IN1(n10375), .IN2(n10376), .Q(n10373) );
  AO221X1 U2747 ( .IN1(\U611/DATA1_3 ), .IN2(n14375), .IN3(\U616/DATA1_3 ), 
        .IN4(n9447), .IN5(n10377), .Q(n10376) );
  AO22X1 U2748 ( .IN1(\U586/DATA1_3 ), .IN2(n14193), .IN3(\U616/DATA2_3 ), 
        .IN4(n14361), .Q(n10377) );
  AO221X1 U2749 ( .IN1(\U591/DATA1_3 ), .IN2(n9451), .IN3(\U606/DATA1_3 ), 
        .IN4(n14334), .IN5(n10378), .Q(n10375) );
  AO22X1 U2750 ( .IN1(\U596/DATA1_3 ), .IN2(n9454), .IN3(\U601/DATA1_3 ), 
        .IN4(n14323), .Q(n10378) );
  AO21X1 U2751 ( .IN1(n5956), .IN2(n14244), .IN3(n9542), .Q(n13397) );
  AO22X1 U2753 ( .IN1(\U571/DATA1_2 ), .IN2(n14258), .IN3(\U581/DATA1_2 ), 
        .IN4(n14394), .Q(n10380) );
  OR2X1 U2754 ( .IN1(n10381), .IN2(n10382), .Q(n10379) );
  AO221X1 U2755 ( .IN1(\U611/DATA1_2 ), .IN2(n9446), .IN3(\U616/DATA1_2 ), 
        .IN4(n14374), .IN5(n10383), .Q(n10382) );
  AO22X1 U2756 ( .IN1(\U586/DATA1_2 ), .IN2(n14257), .IN3(\U616/DATA2_2 ), 
        .IN4(n9450), .Q(n10383) );
  AO221X1 U2757 ( .IN1(\U591/DATA1_2 ), .IN2(n9451), .IN3(\U606/DATA1_2 ), 
        .IN4(n14342), .IN5(n10384), .Q(n10381) );
  AO22X1 U2758 ( .IN1(\U596/DATA1_2 ), .IN2(n14324), .IN3(\U601/DATA1_2 ), 
        .IN4(n9455), .Q(n10384) );
  AO21X1 U2759 ( .IN1(n5955), .IN2(n14239), .IN3(n9544), .Q(n13398) );
  AO22X1 U2761 ( .IN1(\U571/DATA1_1 ), .IN2(n14258), .IN3(\U581/DATA1_1 ), 
        .IN4(n14394), .Q(n10386) );
  OR2X1 U2762 ( .IN1(n10387), .IN2(n10388), .Q(n10385) );
  AO221X1 U2763 ( .IN1(\U611/DATA1_1 ), .IN2(n9446), .IN3(\U616/DATA1_1 ), 
        .IN4(n9447), .IN5(n10389), .Q(n10388) );
  AO22X1 U2764 ( .IN1(\U586/DATA1_1 ), .IN2(n14255), .IN3(\U616/DATA2_1 ), 
        .IN4(n9450), .Q(n10389) );
  AO221X1 U2765 ( .IN1(\U591/DATA1_1 ), .IN2(n9451), .IN3(\U606/DATA1_1 ), 
        .IN4(n9452), .IN5(n10390), .Q(n10387) );
  AO22X1 U2766 ( .IN1(\U596/DATA1_1 ), .IN2(n9454), .IN3(\U601/DATA1_1 ), 
        .IN4(n9455), .Q(n10390) );
  AO22X1 U2769 ( .IN1(\U581/DATA1_0 ), .IN2(n14394), .IN3(\U576/DATA1_0 ), 
        .IN4(n9440), .Q(n10392) );
  OR2X1 U2773 ( .IN1(n10394), .IN2(n10395), .Q(n10391) );
  AO221X1 U2774 ( .IN1(\U611/DATA1_0 ), .IN2(n9446), .IN3(\U616/DATA1_0 ), 
        .IN4(n14364), .IN5(n10396), .Q(n10395) );
  AO22X1 U2775 ( .IN1(\U586/DATA1_0 ), .IN2(n14256), .IN3(\U616/DATA2_0 ), 
        .IN4(n9450), .Q(n10396) );
  NOR3X0 U2776 ( .IN1(n10397), .IN2(n12837), .IN3(n13537), .QN(n9447) );
  AO221X1 U2778 ( .IN1(\U591/DATA1_0 ), .IN2(n9451), .IN3(\U606/DATA1_0 ), 
        .IN4(n14334), .IN5(n10399), .Q(n10394) );
  AO22X1 U2779 ( .IN1(\U596/DATA1_0 ), .IN2(n14325), .IN3(\U601/DATA1_0 ), 
        .IN4(n9455), .Q(n10399) );
  NOR3X0 U2780 ( .IN1(n10400), .IN2(n12834), .IN3(n13698), .QN(n9455) );
  AND3X1 U2786 ( .IN1(n14915), .IN2(n10404), .IN3(n12831), .Q(n9441) );
  NAND4X0 U2788 ( .IN1(n12831), .IN2(n9450), .IN3(n14915), .IN4(n13715), .QN(
        n10404) );
  NOR3X0 U2791 ( .IN1(n13674), .IN2(n10397), .IN3(n13537), .QN(n9450) );
  NAND3X0 U2795 ( .IN1(n12834), .IN2(n14913), .IN3(n12833), .QN(n10402) );
  AO22X1 U2822 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/B[1] ), 
        .IN2(\fmul_0_0_0_0_9/sigprod [8]), .IN3(\fmul_0_0_0_0_9/sigprod [7]), 
        .IN4(\add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/B[0] ), .Q(
        \fmul_0_0_0_0_9/sigprodext [9]) );
  AO22X1 U2823 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/B[1] ), 
        .IN2(\fmul_0_0_0_0_9/sigprod [7]), .IN3(\fmul_0_0_0_0_9/sigprod [6]), 
        .IN4(\add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/B[0] ), .Q(
        \fmul_0_0_0_0_9/sigprodext [8]) );
  AO22X1 U2824 ( .IN1(\fmul_0_0_0_0_9/sigprod [6]), .IN2(
        \add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/B[1] ), .IN3(
        \fmul_0_0_0_0_9/sigprod [5]), .IN4(
        \add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/B[0] ), .Q(
        \fmul_0_0_0_0_9/sigprodext [7]) );
  AO22X1 U2825 ( .IN1(\fmul_0_0_0_0_9/sigprod [5]), .IN2(
        \add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/B[1] ), .IN3(
        \fmul_0_0_0_0_9/sigprod [4]), .IN4(
        \add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/B[0] ), .Q(
        \fmul_0_0_0_0_9/sigprodext [6]) );
  XOR2X1 U2826 ( .IN1(n11648), .IN2(n11649), .Q(\fmul_0_0_0_0_9/sign ) );
  NAND3X0 U2828 ( .IN1(n10424), .IN2(
        \add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/B[0] ), .IN3(
        \fmul_0_0_0_0_9/sigprod [3]), .QN(n10423) );
  OAI21X1 U2830 ( .IN1(\fmul_0_0_0_0_9/sigprod [3]), .IN2(n10425), .IN3(
        \fmul_0_0_0_0_9/sigprod [4]), .QN(n10422) );
  OA21X1 U2831 ( .IN1(n10424), .IN2(\fmul_0_0_0_0_9/sigprod [5]), .IN3(
        \add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/B[1] ), .Q(n10425) );
  OR3X1 U2832 ( .IN1(\fmul_0_0_0_0_9/sigprod [2]), .IN2(
        \fmul_0_0_0_0_9/sigprod [1]), .IN3(\fmul_0_0_0_0_9/sigprod [0]), .Q(
        n10424) );
  AO22X1 U2833 ( .IN1(n13896), .IN2(n13606), .IN3(n10426), .IN4(
        \fmul_0_0_0_0_9/exc [1]), .Q(\fmul_0_0_0_0_9/exc [0]) );
  OA21X1 U2835 ( .IN1(n12788), .IN2(n13764), .IN3(n10427), .Q(n10426) );
  NAND3X0 U2836 ( .IN1(n10428), .IN2(n13764), .IN3(n12788), .QN(n10427) );
  XOR2X1 U2837 ( .IN1(n11650), .IN2(n11651), .Q(n10428) );
  AO22X1 U2841 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/B[1] ), 
        .IN2(\fmul_0_0_0_0_8/sigprod [8]), .IN3(\fmul_0_0_0_0_8/sigprod [7]), 
        .IN4(\add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/B[0] ), .Q(
        \fmul_0_0_0_0_8/sigprodext [9]) );
  AO22X1 U2842 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/B[1] ), 
        .IN2(\fmul_0_0_0_0_8/sigprod [7]), .IN3(\fmul_0_0_0_0_8/sigprod [6]), 
        .IN4(\add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/B[0] ), .Q(
        \fmul_0_0_0_0_8/sigprodext [8]) );
  AO22X1 U2843 ( .IN1(\fmul_0_0_0_0_8/sigprod [6]), .IN2(
        \add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/B[1] ), .IN3(
        \fmul_0_0_0_0_8/sigprod [5]), .IN4(
        \add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/B[0] ), .Q(
        \fmul_0_0_0_0_8/sigprodext [7]) );
  AO22X1 U2844 ( .IN1(\fmul_0_0_0_0_8/sigprod [5]), .IN2(
        \add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/B[1] ), .IN3(
        \fmul_0_0_0_0_8/sigprod [4]), .IN4(
        \add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/B[0] ), .Q(
        \fmul_0_0_0_0_8/sigprodext [6]) );
  XOR2X1 U2845 ( .IN1(n11644), .IN2(n11645), .Q(\fmul_0_0_0_0_8/sign ) );
  NAND3X0 U2847 ( .IN1(n10432), .IN2(
        \add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/B[0] ), .IN3(
        \fmul_0_0_0_0_8/sigprod [3]), .QN(n10431) );
  OAI21X1 U2849 ( .IN1(\fmul_0_0_0_0_8/sigprod [3]), .IN2(n10433), .IN3(
        \fmul_0_0_0_0_8/sigprod [4]), .QN(n10430) );
  OA21X1 U2850 ( .IN1(n10432), .IN2(\fmul_0_0_0_0_8/sigprod [5]), .IN3(
        \add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/B[1] ), .Q(n10433) );
  OR3X1 U2851 ( .IN1(\fmul_0_0_0_0_8/sigprod [2]), .IN2(
        \fmul_0_0_0_0_8/sigprod [1]), .IN3(\fmul_0_0_0_0_8/sigprod [0]), .Q(
        n10432) );
  AO22X1 U2852 ( .IN1(n13895), .IN2(n13605), .IN3(n10434), .IN4(
        \fmul_0_0_0_0_8/exc [1]), .Q(\fmul_0_0_0_0_8/exc [0]) );
  OA21X1 U2854 ( .IN1(n12778), .IN2(n13763), .IN3(n10435), .Q(n10434) );
  NAND3X0 U2855 ( .IN1(n10436), .IN2(n13763), .IN3(n12778), .QN(n10435) );
  XOR2X1 U2856 ( .IN1(n11646), .IN2(n11647), .Q(n10436) );
  AO22X1 U2860 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/B[1] ), 
        .IN2(\fmul_0_0_0_0_7/sigprod [8]), .IN3(\fmul_0_0_0_0_7/sigprod [7]), 
        .IN4(\add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/B[0] ), .Q(
        \fmul_0_0_0_0_7/sigprodext [9]) );
  AO22X1 U2861 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/B[1] ), 
        .IN2(\fmul_0_0_0_0_7/sigprod [7]), .IN3(\fmul_0_0_0_0_7/sigprod [6]), 
        .IN4(\add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/B[0] ), .Q(
        \fmul_0_0_0_0_7/sigprodext [8]) );
  AO22X1 U2862 ( .IN1(\fmul_0_0_0_0_7/sigprod [6]), .IN2(
        \add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/B[1] ), .IN3(
        \fmul_0_0_0_0_7/sigprod [5]), .IN4(
        \add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/B[0] ), .Q(
        \fmul_0_0_0_0_7/sigprodext [7]) );
  AO22X1 U2863 ( .IN1(\fmul_0_0_0_0_7/sigprod [5]), .IN2(
        \add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/B[1] ), .IN3(
        \fmul_0_0_0_0_7/sigprod [4]), .IN4(
        \add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/B[0] ), .Q(
        \fmul_0_0_0_0_7/sigprodext [6]) );
  XOR2X1 U2864 ( .IN1(n11640), .IN2(n11641), .Q(\fmul_0_0_0_0_7/sign ) );
  NAND3X0 U2866 ( .IN1(n10440), .IN2(
        \add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/B[0] ), .IN3(
        \fmul_0_0_0_0_7/sigprod [3]), .QN(n10439) );
  OAI21X1 U2868 ( .IN1(\fmul_0_0_0_0_7/sigprod [3]), .IN2(n10441), .IN3(
        \fmul_0_0_0_0_7/sigprod [4]), .QN(n10438) );
  OA21X1 U2869 ( .IN1(n10440), .IN2(\fmul_0_0_0_0_7/sigprod [5]), .IN3(
        \add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/B[1] ), .Q(n10441) );
  OR3X1 U2870 ( .IN1(\fmul_0_0_0_0_7/sigprod [2]), .IN2(
        \fmul_0_0_0_0_7/sigprod [1]), .IN3(\fmul_0_0_0_0_7/sigprod [0]), .Q(
        n10440) );
  AO22X1 U2871 ( .IN1(n13615), .IN2(n13905), .IN3(n10442), .IN4(
        \fmul_0_0_0_0_7/exc [1]), .Q(\fmul_0_0_0_0_7/exc [0]) );
  OA21X1 U2873 ( .IN1(n12768), .IN2(n13762), .IN3(n10443), .Q(n10442) );
  NAND3X0 U2874 ( .IN1(n10444), .IN2(n13762), .IN3(n12768), .QN(n10443) );
  XOR2X1 U2875 ( .IN1(n11642), .IN2(n11643), .Q(n10444) );
  AO22X1 U2879 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/B[1] ), 
        .IN2(\fmul_0_0_0_0_6/sigprod [8]), .IN3(\fmul_0_0_0_0_6/sigprod [7]), 
        .IN4(\add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/B[0] ), .Q(
        \fmul_0_0_0_0_6/sigprodext [9]) );
  AO22X1 U2880 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/B[1] ), 
        .IN2(\fmul_0_0_0_0_6/sigprod [7]), .IN3(\fmul_0_0_0_0_6/sigprod [6]), 
        .IN4(\add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/B[0] ), .Q(
        \fmul_0_0_0_0_6/sigprodext [8]) );
  AO22X1 U2881 ( .IN1(\fmul_0_0_0_0_6/sigprod [6]), .IN2(
        \add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/B[1] ), .IN3(
        \fmul_0_0_0_0_6/sigprod [5]), .IN4(
        \add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/B[0] ), .Q(
        \fmul_0_0_0_0_6/sigprodext [7]) );
  AO22X1 U2882 ( .IN1(\fmul_0_0_0_0_6/sigprod [5]), .IN2(
        \add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/B[1] ), .IN3(
        \fmul_0_0_0_0_6/sigprod [4]), .IN4(
        \add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/B[0] ), .Q(
        \fmul_0_0_0_0_6/sigprodext [6]) );
  XOR2X1 U2883 ( .IN1(n11636), .IN2(n11637), .Q(\fmul_0_0_0_0_6/sign ) );
  NAND3X0 U2885 ( .IN1(n10448), .IN2(
        \add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/B[0] ), .IN3(
        \fmul_0_0_0_0_6/sigprod [3]), .QN(n10447) );
  OAI21X1 U2887 ( .IN1(\fmul_0_0_0_0_6/sigprod [3]), .IN2(n10449), .IN3(
        \fmul_0_0_0_0_6/sigprod [4]), .QN(n10446) );
  OA21X1 U2888 ( .IN1(n10448), .IN2(\fmul_0_0_0_0_6/sigprod [5]), .IN3(
        \add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/B[1] ), .Q(n10449) );
  OR3X1 U2889 ( .IN1(\fmul_0_0_0_0_6/sigprod [2]), .IN2(
        \fmul_0_0_0_0_6/sigprod [1]), .IN3(\fmul_0_0_0_0_6/sigprod [0]), .Q(
        n10448) );
  AO22X1 U2890 ( .IN1(n13614), .IN2(n13904), .IN3(n10450), .IN4(
        \fmul_0_0_0_0_6/exc [1]), .Q(\fmul_0_0_0_0_6/exc [0]) );
  OA21X1 U2892 ( .IN1(n12750), .IN2(n13761), .IN3(n10451), .Q(n10450) );
  NAND3X0 U2893 ( .IN1(n10452), .IN2(n13761), .IN3(n12750), .QN(n10451) );
  XOR2X1 U2894 ( .IN1(n11638), .IN2(n11639), .Q(n10452) );
  AO22X1 U2898 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/B[1] ), 
        .IN2(\fmul_0_0_0_0_5/sigprod [8]), .IN3(\fmul_0_0_0_0_5/sigprod [7]), 
        .IN4(\add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/B[0] ), .Q(
        \fmul_0_0_0_0_5/sigprodext [9]) );
  AO22X1 U2899 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/B[1] ), 
        .IN2(\fmul_0_0_0_0_5/sigprod [7]), .IN3(\fmul_0_0_0_0_5/sigprod [6]), 
        .IN4(\add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/B[0] ), .Q(
        \fmul_0_0_0_0_5/sigprodext [8]) );
  AO22X1 U2900 ( .IN1(\fmul_0_0_0_0_5/sigprod [6]), .IN2(
        \add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/B[1] ), .IN3(
        \fmul_0_0_0_0_5/sigprod [5]), .IN4(
        \add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/B[0] ), .Q(
        \fmul_0_0_0_0_5/sigprodext [7]) );
  AO22X1 U2901 ( .IN1(\fmul_0_0_0_0_5/sigprod [5]), .IN2(
        \add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/B[1] ), .IN3(
        \fmul_0_0_0_0_5/sigprod [4]), .IN4(
        \add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/B[0] ), .Q(
        \fmul_0_0_0_0_5/sigprodext [6]) );
  XOR2X1 U2902 ( .IN1(n11632), .IN2(n11633), .Q(\fmul_0_0_0_0_5/sign ) );
  NAND3X0 U2904 ( .IN1(n10456), .IN2(
        \add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/B[0] ), .IN3(
        \fmul_0_0_0_0_5/sigprod [3]), .QN(n10455) );
  OAI21X1 U2906 ( .IN1(\fmul_0_0_0_0_5/sigprod [3]), .IN2(n10457), .IN3(
        \fmul_0_0_0_0_5/sigprod [4]), .QN(n10454) );
  OA21X1 U2907 ( .IN1(n10456), .IN2(\fmul_0_0_0_0_5/sigprod [5]), .IN3(
        \add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/B[1] ), .Q(n10457) );
  OR3X1 U2908 ( .IN1(\fmul_0_0_0_0_5/sigprod [2]), .IN2(
        \fmul_0_0_0_0_5/sigprod [1]), .IN3(\fmul_0_0_0_0_5/sigprod [0]), .Q(
        n10456) );
  AO22X1 U2909 ( .IN1(n13613), .IN2(n13903), .IN3(n10458), .IN4(
        \fmul_0_0_0_0_5/exc [1]), .Q(\fmul_0_0_0_0_5/exc [0]) );
  OA21X1 U2911 ( .IN1(n12748), .IN2(n13760), .IN3(n10459), .Q(n10458) );
  NAND3X0 U2912 ( .IN1(n10460), .IN2(n13760), .IN3(n12748), .QN(n10459) );
  XOR2X1 U2913 ( .IN1(n11634), .IN2(n11635), .Q(n10460) );
  AO22X1 U2917 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/B[1] ), 
        .IN2(\fmul_0_0_0_0_4/sigprod [8]), .IN3(\fmul_0_0_0_0_4/sigprod [7]), 
        .IN4(\add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/B[0] ), .Q(
        \fmul_0_0_0_0_4/sigprodext [9]) );
  AO22X1 U2918 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/B[1] ), 
        .IN2(\fmul_0_0_0_0_4/sigprod [7]), .IN3(\fmul_0_0_0_0_4/sigprod [6]), 
        .IN4(\add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/B[0] ), .Q(
        \fmul_0_0_0_0_4/sigprodext [8]) );
  AO22X1 U2919 ( .IN1(\fmul_0_0_0_0_4/sigprod [6]), .IN2(
        \add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/B[1] ), .IN3(
        \fmul_0_0_0_0_4/sigprod [5]), .IN4(
        \add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/B[0] ), .Q(
        \fmul_0_0_0_0_4/sigprodext [7]) );
  AO22X1 U2920 ( .IN1(\fmul_0_0_0_0_4/sigprod [5]), .IN2(
        \add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/B[1] ), .IN3(
        \fmul_0_0_0_0_4/sigprod [4]), .IN4(
        \add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/B[0] ), .Q(
        \fmul_0_0_0_0_4/sigprodext [6]) );
  XOR2X1 U2921 ( .IN1(n11628), .IN2(n11629), .Q(\fmul_0_0_0_0_4/sign ) );
  NAND3X0 U2923 ( .IN1(n10464), .IN2(
        \add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/B[0] ), .IN3(
        \fmul_0_0_0_0_4/sigprod [3]), .QN(n10463) );
  OAI21X1 U2925 ( .IN1(\fmul_0_0_0_0_4/sigprod [3]), .IN2(n10465), .IN3(
        \fmul_0_0_0_0_4/sigprod [4]), .QN(n10462) );
  OA21X1 U2926 ( .IN1(n10464), .IN2(\fmul_0_0_0_0_4/sigprod [5]), .IN3(
        \add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/B[1] ), .Q(n10465) );
  OR3X1 U2927 ( .IN1(\fmul_0_0_0_0_4/sigprod [2]), .IN2(
        \fmul_0_0_0_0_4/sigprod [1]), .IN3(\fmul_0_0_0_0_4/sigprod [0]), .Q(
        n10464) );
  AO22X1 U2928 ( .IN1(n13612), .IN2(n13902), .IN3(n10466), .IN4(
        \fmul_0_0_0_0_4/exc [1]), .Q(\fmul_0_0_0_0_4/exc [0]) );
  OA21X1 U2930 ( .IN1(n12730), .IN2(n13759), .IN3(n10467), .Q(n10466) );
  NAND3X0 U2931 ( .IN1(n10468), .IN2(n13759), .IN3(n12730), .QN(n10467) );
  XOR2X1 U2932 ( .IN1(n11630), .IN2(n11631), .Q(n10468) );
  AO22X1 U2936 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/B[1] ), 
        .IN2(\fmul_0_0_0_0_3/sigprod [8]), .IN3(\fmul_0_0_0_0_3/sigprod [7]), 
        .IN4(\add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/B[0] ), .Q(
        \fmul_0_0_0_0_3/sigprodext [9]) );
  AO22X1 U2937 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/B[1] ), 
        .IN2(\fmul_0_0_0_0_3/sigprod [7]), .IN3(\fmul_0_0_0_0_3/sigprod [6]), 
        .IN4(\add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/B[0] ), .Q(
        \fmul_0_0_0_0_3/sigprodext [8]) );
  AO22X1 U2938 ( .IN1(\fmul_0_0_0_0_3/sigprod [6]), .IN2(
        \add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/B[1] ), .IN3(
        \fmul_0_0_0_0_3/sigprod [5]), .IN4(
        \add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/B[0] ), .Q(
        \fmul_0_0_0_0_3/sigprodext [7]) );
  AO22X1 U2939 ( .IN1(\fmul_0_0_0_0_3/sigprod [5]), .IN2(
        \add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/B[1] ), .IN3(
        \fmul_0_0_0_0_3/sigprod [4]), .IN4(
        \add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/B[0] ), .Q(
        \fmul_0_0_0_0_3/sigprodext [6]) );
  XOR2X1 U2940 ( .IN1(n11624), .IN2(n11625), .Q(\fmul_0_0_0_0_3/sign ) );
  NAND3X0 U2942 ( .IN1(n10472), .IN2(
        \add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/B[0] ), .IN3(
        \fmul_0_0_0_0_3/sigprod [3]), .QN(n10471) );
  OAI21X1 U2944 ( .IN1(\fmul_0_0_0_0_3/sigprod [3]), .IN2(n10473), .IN3(
        \fmul_0_0_0_0_3/sigprod [4]), .QN(n10470) );
  OA21X1 U2945 ( .IN1(n10472), .IN2(\fmul_0_0_0_0_3/sigprod [5]), .IN3(
        \add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/B[1] ), .Q(n10473) );
  OR3X1 U2946 ( .IN1(\fmul_0_0_0_0_3/sigprod [2]), .IN2(
        \fmul_0_0_0_0_3/sigprod [1]), .IN3(\fmul_0_0_0_0_3/sigprod [0]), .Q(
        n10472) );
  AO22X1 U2947 ( .IN1(n13611), .IN2(n13901), .IN3(n10474), .IN4(
        \fmul_0_0_0_0_3/exc [1]), .Q(\fmul_0_0_0_0_3/exc [0]) );
  OA21X1 U2949 ( .IN1(n12728), .IN2(n13758), .IN3(n10475), .Q(n10474) );
  NAND3X0 U2950 ( .IN1(n10476), .IN2(n13758), .IN3(n12728), .QN(n10475) );
  XOR2X1 U2951 ( .IN1(n11626), .IN2(n11627), .Q(n10476) );
  AO22X1 U2955 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/B[1] ), 
        .IN2(\fmul_0_0_0_0_2/sigprod [8]), .IN3(\fmul_0_0_0_0_2/sigprod [7]), 
        .IN4(\add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/B[0] ), .Q(
        \fmul_0_0_0_0_2/sigprodext [9]) );
  AO22X1 U2956 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/B[1] ), 
        .IN2(\fmul_0_0_0_0_2/sigprod [7]), .IN3(\fmul_0_0_0_0_2/sigprod [6]), 
        .IN4(\add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/B[0] ), .Q(
        \fmul_0_0_0_0_2/sigprodext [8]) );
  AO22X1 U2957 ( .IN1(\fmul_0_0_0_0_2/sigprod [6]), .IN2(
        \add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/B[1] ), .IN3(
        \fmul_0_0_0_0_2/sigprod [5]), .IN4(
        \add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/B[0] ), .Q(
        \fmul_0_0_0_0_2/sigprodext [7]) );
  AO22X1 U2958 ( .IN1(\fmul_0_0_0_0_2/sigprod [5]), .IN2(
        \add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/B[1] ), .IN3(
        \fmul_0_0_0_0_2/sigprod [4]), .IN4(
        \add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/B[0] ), .Q(
        \fmul_0_0_0_0_2/sigprodext [6]) );
  XOR2X1 U2959 ( .IN1(n11620), .IN2(n11621), .Q(\fmul_0_0_0_0_2/sign ) );
  NAND3X0 U2961 ( .IN1(n10480), .IN2(
        \add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/B[0] ), .IN3(
        \fmul_0_0_0_0_2/sigprod [3]), .QN(n10479) );
  OAI21X1 U2963 ( .IN1(\fmul_0_0_0_0_2/sigprod [3]), .IN2(n10481), .IN3(
        \fmul_0_0_0_0_2/sigprod [4]), .QN(n10478) );
  OA21X1 U2964 ( .IN1(n10480), .IN2(\fmul_0_0_0_0_2/sigprod [5]), .IN3(
        \add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/B[1] ), .Q(n10481) );
  OR3X1 U2965 ( .IN1(\fmul_0_0_0_0_2/sigprod [2]), .IN2(
        \fmul_0_0_0_0_2/sigprod [1]), .IN3(\fmul_0_0_0_0_2/sigprod [0]), .Q(
        n10480) );
  AO22X1 U2966 ( .IN1(n13610), .IN2(n13900), .IN3(n10482), .IN4(
        \fmul_0_0_0_0_2/exc [1]), .Q(\fmul_0_0_0_0_2/exc [0]) );
  OA21X1 U2968 ( .IN1(n12710), .IN2(n13757), .IN3(n10483), .Q(n10482) );
  NAND3X0 U2969 ( .IN1(n10484), .IN2(n13757), .IN3(n12710), .QN(n10483) );
  XOR2X1 U2970 ( .IN1(n11622), .IN2(n11623), .Q(n10484) );
  AOI22X1 U2975 ( .IN1(n10487), .IN2(n10488), .IN3(n14920), .IN4(n10489), .QN(
        n10486) );
  NOR3X0 U2976 ( .IN1(n10490), .IN2(n10491), .IN3(n10492), .QN(n10485) );
  AO221X1 U2978 ( .IN1(n10493), .IN2(n13618), .IN3(n10488), .IN4(n14920), 
        .IN5(\fmul_0_0_0_0_10/U8/Z_5 ), .Q(n10490) );
  XOR2X1 U2979 ( .IN1(n10494), .IN2(n10495), .Q(n10488) );
  XOR2X1 U2981 ( .IN1(n11652), .IN2(n11653), .Q(\fmul_0_0_0_0_10/n137 ) );
  AO22X1 U2982 ( .IN1(n13897), .IN2(n13607), .IN3(n10496), .IN4(
        \fmul_0_0_0_0_10/U9/Z_1 ), .Q(\fmul_0_0_0_0_10/U9/Z_0 ) );
  OA21X1 U2984 ( .IN1(n12816), .IN2(n13765), .IN3(n10497), .Q(n10496) );
  NAND3X0 U2985 ( .IN1(n10498), .IN2(n13765), .IN3(n12816), .QN(n10497) );
  XOR2X1 U2986 ( .IN1(n11654), .IN2(n11655), .Q(n10498) );
  AO22X1 U2990 ( .IN1(n10499), .IN2(n10487), .IN3(n10500), .IN4(n14922), .Q(
        \fmul_0_0_0_0_10/U8/Z_8 ) );
  AO22X1 U2993 ( .IN1(n10505), .IN2(n10487), .IN3(n10499), .IN4(n14920), .Q(
        \fmul_0_0_0_0_10/U8/Z_7 ) );
  AO222X1 U2994 ( .IN1(n10506), .IN2(n10507), .IN3(n14923), .IN4(n14921), 
        .IN5(n10502), .IN6(n10509), .Q(n10499) );
  AO22X1 U2996 ( .IN1(n10511), .IN2(n10487), .IN3(n10505), .IN4(n14920), .Q(
        \fmul_0_0_0_0_10/U8/Z_6 ) );
  XOR3X1 U2997 ( .IN1(n10512), .IN2(n10513), .IN3(n10514), .Q(n10505) );
  AO22X1 U2998 ( .IN1(n10511), .IN2(n14920), .IN3(n10489), .IN4(n10487), .Q(
        \fmul_0_0_0_0_10/U8/Z_5 ) );
  XOR3X1 U2999 ( .IN1(n10515), .IN2(n10516), .IN3(n10517), .Q(n10489) );
  OA21X1 U3001 ( .IN1(n14921), .IN2(n10502), .IN3(n10503), .Q(n10487) );
  AOI21X1 U3002 ( .IN1(n10518), .IN2(n10519), .IN3(n14925), .QN(n10503) );
  AO21X1 U3006 ( .IN1(n10521), .IN2(n10522), .IN3(n10523), .Q(n10510) );
  AO22X1 U3007 ( .IN1(n10512), .IN2(n10513), .IN3(n10524), .IN4(n10514), .Q(
        n10507) );
  AO22X1 U3008 ( .IN1(n10525), .IN2(n10526), .IN3(n10527), .IN4(n10528), .Q(
        n10514) );
  OR2X1 U3009 ( .IN1(n10526), .IN2(n10525), .Q(n10528) );
  OR2X1 U3010 ( .IN1(n10513), .IN2(n10512), .Q(n10524) );
  AO22X1 U3011 ( .IN1(n10529), .IN2(n10530), .IN3(n10531), .IN4(n10532), .Q(
        n10513) );
  OR2X1 U3012 ( .IN1(n10529), .IN2(n10530), .Q(n10532) );
  XNOR3X1 U3013 ( .IN1(n10521), .IN2(n10523), .IN3(n10522), .Q(n10512) );
  AO22X1 U3014 ( .IN1(n10533), .IN2(n10534), .IN3(n12821), .IN4(n10535), .Q(
        n10522) );
  OR2X1 U3015 ( .IN1(n10534), .IN2(n10533), .Q(n10535) );
  AO222X1 U3016 ( .IN1(n10536), .IN2(n14925), .IN3(n12824), .IN4(n10537), 
        .IN5(n10538), .IN6(n10539), .Q(n10523) );
  XOR2X1 U3017 ( .IN1(n12820), .IN2(n14925), .Q(n10537) );
  AO222X1 U3021 ( .IN1(n11924), .IN2(n10541), .IN3(n10542), .IN4(n14924), 
        .IN5(n14925), .IN6(n10519), .Q(n10509) );
  XOR2X1 U3024 ( .IN1(n13499), .IN2(n10519), .Q(n10541) );
  AO21X1 U3025 ( .IN1(n14925), .IN2(n10544), .IN3(n10538), .Q(n10519) );
  XOR3X1 U3029 ( .IN1(n10527), .IN2(n10525), .IN3(n10526), .Q(n10511) );
  AO22X1 U3030 ( .IN1(n10515), .IN2(n10516), .IN3(n10545), .IN4(n10517), .Q(
        n10526) );
  AO22X1 U3031 ( .IN1(n10495), .IN2(n10494), .IN3(n14926), .IN4(n14927), .Q(
        n10517) );
  NAND3X0 U3035 ( .IN1(n13620), .IN2(n13498), .IN3(n10550), .QN(n10548) );
  AO22X1 U3037 ( .IN1(n10492), .IN2(n13619), .IN3(n10552), .IN4(n10553), .Q(
        n10551) );
  OA21X1 U3038 ( .IN1(n13619), .IN2(n10492), .IN3(n13498), .Q(n10552) );
  XNOR2X1 U3039 ( .IN1(n10554), .IN2(n10553), .Q(n10492) );
  XOR3X1 U3043 ( .IN1(n10550), .IN2(n10555), .IN3(n10556), .Q(n10495) );
  OR2X1 U3044 ( .IN1(n10516), .IN2(n10515), .Q(n10545) );
  AO22X1 U3045 ( .IN1(n10555), .IN2(n10556), .IN3(n10550), .IN4(n10557), .Q(
        n10516) );
  OR2X1 U3046 ( .IN1(n10556), .IN2(n10555), .Q(n10557) );
  XNOR2X1 U3048 ( .IN1(n10558), .IN2(n10559), .Q(n10556) );
  XNOR2X1 U3051 ( .IN1(n10560), .IN2(n10561), .Q(n10515) );
  OA21X1 U3053 ( .IN1(n10562), .IN2(n10563), .IN3(n10560), .Q(n10525) );
  XOR3X1 U3054 ( .IN1(n10564), .IN2(n13498), .IN3(n10538), .Q(n10560) );
  AND2X1 U3055 ( .IN1(n10531), .IN2(n13619), .Q(n10563) );
  OA21X1 U3057 ( .IN1(n11924), .IN2(n12825), .IN3(n11923), .Q(n10565) );
  XOR3X1 U3058 ( .IN1(n10531), .IN2(n10530), .IN3(n10529), .Q(n10527) );
  XOR3X1 U3059 ( .IN1(n13629), .IN2(n10534), .IN3(n10533), .Q(n10529) );
  XNOR2X1 U3060 ( .IN1(n13620), .IN2(n10540), .Q(n10533) );
  AO22X1 U3067 ( .IN1(n10564), .IN2(n10538), .IN3(n10566), .IN4(n13498), .Q(
        n10530) );
  OR2X1 U3069 ( .IN1(n10564), .IN2(n10538), .Q(n10566) );
  AO22X1 U3076 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/B[1] ), 
        .IN2(\fmul_0_0_0_0_1/sigprod [8]), .IN3(\fmul_0_0_0_0_1/sigprod [7]), 
        .IN4(\add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/B[0] ), .Q(
        \fmul_0_0_0_0_1/sigprodext [9]) );
  AO22X1 U3077 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/B[1] ), 
        .IN2(\fmul_0_0_0_0_1/sigprod [7]), .IN3(\fmul_0_0_0_0_1/sigprod [6]), 
        .IN4(\add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/B[0] ), .Q(
        \fmul_0_0_0_0_1/sigprodext [8]) );
  AO22X1 U3078 ( .IN1(\fmul_0_0_0_0_1/sigprod [6]), .IN2(
        \add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/B[1] ), .IN3(
        \fmul_0_0_0_0_1/sigprod [5]), .IN4(
        \add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/B[0] ), .Q(
        \fmul_0_0_0_0_1/sigprodext [7]) );
  AO22X1 U3079 ( .IN1(\fmul_0_0_0_0_1/sigprod [5]), .IN2(
        \add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/B[1] ), .IN3(
        \fmul_0_0_0_0_1/sigprod [4]), .IN4(
        \add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/B[0] ), .Q(
        \fmul_0_0_0_0_1/sigprodext [6]) );
  XOR2X1 U3080 ( .IN1(n11616), .IN2(n11617), .Q(\fmul_0_0_0_0_1/sign ) );
  NAND3X0 U3082 ( .IN1(n10570), .IN2(
        \add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/B[0] ), .IN3(
        \fmul_0_0_0_0_1/sigprod [3]), .QN(n10569) );
  OAI21X1 U3084 ( .IN1(\fmul_0_0_0_0_1/sigprod [3]), .IN2(n10571), .IN3(
        \fmul_0_0_0_0_1/sigprod [4]), .QN(n10568) );
  OA21X1 U3085 ( .IN1(n10570), .IN2(\fmul_0_0_0_0_1/sigprod [5]), .IN3(
        \add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/B[1] ), .Q(n10571) );
  OR3X1 U3086 ( .IN1(\fmul_0_0_0_0_1/sigprod [2]), .IN2(
        \fmul_0_0_0_0_1/sigprod [1]), .IN3(\fmul_0_0_0_0_1/sigprod [0]), .Q(
        n10570) );
  AO22X1 U3087 ( .IN1(n13609), .IN2(n13899), .IN3(n10572), .IN4(
        \fmul_0_0_0_0_1/exc [1]), .Q(\fmul_0_0_0_0_1/exc [0]) );
  OA21X1 U3089 ( .IN1(n12708), .IN2(n13756), .IN3(n10573), .Q(n10572) );
  NAND3X0 U3090 ( .IN1(n10574), .IN2(n13756), .IN3(n12708), .QN(n10573) );
  XOR2X1 U3091 ( .IN1(n11618), .IN2(n11619), .Q(n10574) );
  AO22X1 U3095 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/B[1] ), 
        .IN2(\fmul_0_0_0_0_0/sigprod [8]), .IN3(\fmul_0_0_0_0_0/sigprod [7]), 
        .IN4(\add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/B[0] ), .Q(
        \fmul_0_0_0_0_0/sigprodext [9]) );
  AO22X1 U3096 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/B[1] ), 
        .IN2(\fmul_0_0_0_0_0/sigprod [7]), .IN3(\fmul_0_0_0_0_0/sigprod [6]), 
        .IN4(\add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/B[0] ), .Q(
        \fmul_0_0_0_0_0/sigprodext [8]) );
  AO22X1 U3097 ( .IN1(\fmul_0_0_0_0_0/sigprod [6]), .IN2(
        \add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/B[1] ), .IN3(
        \fmul_0_0_0_0_0/sigprod [5]), .IN4(
        \add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/B[0] ), .Q(
        \fmul_0_0_0_0_0/sigprodext [7]) );
  XOR2X1 U3098 ( .IN1(n11612), .IN2(n11613), .Q(\fmul_0_0_0_0_0/sign ) );
  AOI22X1 U3100 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/B[0] ), 
        .IN2(\fmul_0_0_0_0_0/sigprod [3]), .IN3(
        \add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/B[1] ), .IN4(
        \fmul_0_0_0_0_0/sigprod [4]), .QN(n10577) );
  AO21X1 U3102 ( .IN1(\fmul_0_0_0_0_0/sigprod [3]), .IN2(
        \add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/B[1] ), .IN3(
        \fmul_0_0_0_0_0/sigprodext [6]), .Q(n10578) );
  AO22X1 U3103 ( .IN1(\fmul_0_0_0_0_0/sigprod [5]), .IN2(
        \add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/B[1] ), .IN3(
        \fmul_0_0_0_0_0/sigprod [4]), .IN4(
        \add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/B[0] ), .Q(
        \fmul_0_0_0_0_0/sigprodext [6]) );
  AO22X1 U3105 ( .IN1(n13608), .IN2(n13898), .IN3(n10579), .IN4(
        \fmul_0_0_0_0_0/exc [1]), .Q(\fmul_0_0_0_0_0/exc [0]) );
  OA21X1 U3107 ( .IN1(n12690), .IN2(n13755), .IN3(n10580), .Q(n10579) );
  NAND3X0 U3108 ( .IN1(n10581), .IN2(n13755), .IN3(n12690), .QN(n10580) );
  XOR2X1 U3109 ( .IN1(n11614), .IN2(n11615), .Q(n10581) );
  NOR3X0 U3113 ( .IN1(n14937), .IN2(n11607), .IN3(n10419), .QN(
        \fadd_0_0_0_0_9/zerofromclose ) );
  NAND3X0 U3115 ( .IN1(n13684), .IN2(n13492), .IN3(n10586), .QN(n10583) );
  NAND3X0 U3116 ( .IN1(n10587), .IN2(n10588), .IN3(n12847), .QN(n10582) );
  AO222X1 U3121 ( .IN1(\fadd_0_0_0_0_9/fracresultfar0 [1]), .IN2(n14891), 
        .IN3(\fadd_0_0_0_0_9/fracresultfar0 [2]), .IN4(n10592), .IN5(
        \fadd_0_0_0_0_9/fracresultfar0 [0]), .IN6(
        \fadd_0_0_0_0_9/add_859/B[1] ), .Q(n10587) );
  AO22X1 U3122 ( .IN1(n10596), .IN2(
        \fadd_0_0_0_0_9/rightshiftercomponent/ps_d1 [1]), .IN3(n10597), .IN4(
        \fadd_0_0_0_0_9/rightshiftercomponent/ps_d1 [2]), .Q(
        \fadd_0_0_0_0_9/rightshiftercomponent/n389_o ) );
  AO22X1 U3125 ( .IN1(n13653), .IN2(\fadd_0_0_0_0_9/exponentresultclose_d1 [5]), .IN3(\fadd_0_0_0_0_9/exponentresultfar1 [5]), .IN4(n12847), .Q(
        \fadd_0_0_0_0_9/resultbeforeround [9]) );
  AO22X1 U3126 ( .IN1(n13653), .IN2(\fadd_0_0_0_0_9/exponentresultclose_d1 [4]), .IN3(\fadd_0_0_0_0_9/exponentresultfar1 [4]), .IN4(n12847), .Q(
        \fadd_0_0_0_0_9/resultbeforeround [8]) );
  AO22X1 U3127 ( .IN1(n13653), .IN2(\fadd_0_0_0_0_9/exponentresultclose_d1 [3]), .IN3(\fadd_0_0_0_0_9/exponentresultfar1 [3]), .IN4(n12847), .Q(
        \fadd_0_0_0_0_9/resultbeforeround [7]) );
  AO22X1 U3128 ( .IN1(n13653), .IN2(\fadd_0_0_0_0_9/exponentresultclose_d1 [2]), .IN3(\fadd_0_0_0_0_9/exponentresultfar1 [2]), .IN4(n12847), .Q(
        \fadd_0_0_0_0_9/resultbeforeround [6]) );
  AO22X1 U3129 ( .IN1(n13653), .IN2(\fadd_0_0_0_0_9/exponentresultclose_d1 [1]), .IN3(\fadd_0_0_0_0_9/exponentresultfar1 [1]), .IN4(n12847), .Q(
        \fadd_0_0_0_0_9/resultbeforeround [5]) );
  AO22X1 U3130 ( .IN1(n13653), .IN2(\fadd_0_0_0_0_9/exponentresultclose_d1 [0]), .IN3(\fadd_0_0_0_0_9/exponentresultfar1 [0]), .IN4(n12847), .Q(
        \fadd_0_0_0_0_9/resultbeforeround [4]) );
  AO222X1 U3131 ( .IN1(n10586), .IN2(\fadd_0_0_0_0_9/norm/level1_d1[4] ), 
        .IN3(n10599), .IN4(n13705), .IN5(n12847), .IN6(n10601), .Q(
        \fadd_0_0_0_0_9/resultbeforeround [3]) );
  AO222X1 U3132 ( .IN1(\fadd_0_0_0_0_9/fracresultfar0 [5]), .IN2(n14891), 
        .IN3(n10592), .IN4(\fadd_0_0_0_0_9/fracresultfar0 [6]), .IN5(
        \fadd_0_0_0_0_9/fracresultfar0 [4]), .IN6(
        \fadd_0_0_0_0_9/add_859/B[1] ), .Q(n10601) );
  AO222X1 U3133 ( .IN1(n10586), .IN2(n13705), .IN3(n10599), .IN4(n13569), 
        .IN5(n12847), .IN6(n10603), .Q(\fadd_0_0_0_0_9/resultbeforeround [2])
         );
  AO222X1 U3134 ( .IN1(\fadd_0_0_0_0_9/fracresultfar0 [4]), .IN2(n14891), 
        .IN3(\fadd_0_0_0_0_9/fracresultfar0 [5]), .IN4(n10592), .IN5(
        \fadd_0_0_0_0_9/add_859/B[1] ), .IN6(
        \fadd_0_0_0_0_9/fracresultfar0 [3]), .Q(n10603) );
  AO222X1 U3136 ( .IN1(n10586), .IN2(n13569), .IN3(n10599), .IN4(n13492), 
        .IN5(n12847), .IN6(n10604), .Q(\fadd_0_0_0_0_9/resultbeforeround [1])
         );
  AO222X1 U3137 ( .IN1(\fadd_0_0_0_0_9/fracresultfar0 [3]), .IN2(n14891), 
        .IN3(\fadd_0_0_0_0_9/fracresultfar0 [4]), .IN4(n10592), .IN5(
        \fadd_0_0_0_0_9/add_859/B[1] ), .IN6(
        \fadd_0_0_0_0_9/fracresultfar0 [2]), .Q(n10604) );
  AO22X1 U3139 ( .IN1(n13653), .IN2(\fadd_0_0_0_0_9/exponentresultclose_d1 [6]), .IN3(\fadd_0_0_0_0_9/exponentresultfar1 [6]), .IN4(n12847), .Q(
        \fadd_0_0_0_0_9/resultbeforeround [10]) );
  AO222X1 U3140 ( .IN1(n10586), .IN2(n13492), .IN3(n10599), .IN4(n13684), 
        .IN5(n12847), .IN6(n10594), .Q(\fadd_0_0_0_0_9/resultbeforeround [0])
         );
  AO222X1 U3141 ( .IN1(\fadd_0_0_0_0_9/fracresultfar0 [2]), .IN2(n14891), 
        .IN3(\fadd_0_0_0_0_9/fracresultfar0 [3]), .IN4(n10592), .IN5(
        \fadd_0_0_0_0_9/fracresultfar0 [1]), .IN6(
        \fadd_0_0_0_0_9/add_859/B[1] ), .Q(n10594) );
  AND2X1 U3148 ( .IN1(n12867), .IN2(n13653), .Q(n10586) );
  OA221X1 U3150 ( .IN1(n10605), .IN2(n10606), .IN3(n10607), .IN4(n10608), 
        .IN5(n10609), .Q(\fadd_0_0_0_0_9/ressign ) );
  XOR2X1 U3151 ( .IN1(n10610), .IN2(n10611), .Q(n10609) );
  OR3X1 U3152 ( .IN1(\fadd_0_0_0_0_9/fracrcloseymx [0]), .IN2(
        \fadd_0_0_0_0_9/fracrcloseymx [1]), .IN3(n10610), .Q(n10608) );
  OR4X1 U3155 ( .IN1(\fadd_0_0_0_0_9/fracrcloseymx [2]), .IN2(
        \fadd_0_0_0_0_9/fracrcloseymx [3]), .IN3(
        \fadd_0_0_0_0_9/fracrcloseymx [4]), .IN4(
        \fadd_0_0_0_0_9/fracrcloseymx [5]), .Q(n10607) );
  OR4X1 U3156 ( .IN1(n10612), .IN2(\fadd_0_0_0_0_9/fracrcloseymx [0]), .IN3(
        \fadd_0_0_0_0_9/fracrclosexmy [1]), .IN4(
        \fadd_0_0_0_0_9/fracrclosexmy [2]), .Q(n10606) );
  AO21X1 U3157 ( .IN1(n10613), .IN2(n10614), .IN3(n14879), .Q(n10612) );
  NAND4X0 U3158 ( .IN1(n10616), .IN2(n10617), .IN3(n14887), .IN4(n14886), .QN(
        n10614) );
  NAND4X0 U3159 ( .IN1(n10620), .IN2(n14312), .IN3(n14889), .IN4(n14888), .QN(
        n10613) );
  AO21X1 U3161 ( .IN1(\fadd_0_0_0_0_9/sub_784/B[1] ), .IN2(n14057), .IN3(
        n10625), .Q(\fadd_0_0_0_0_9/norm/level1 [4]) );
  OAI22X1 U3163 ( .IN1(n14937), .IN2(n11598), .IN3(n10626), .IN4(n11921), .QN(
        \fadd_0_0_0_0_9/norm/level1 [3]) );
  OAI22X1 U3164 ( .IN1(n14937), .IN2(n11597), .IN3(n10626), .IN4(n11922), .QN(
        \fadd_0_0_0_0_9/norm/level1 [2]) );
  NOR3X0 U3169 ( .IN1(n13539), .IN2(n8668), .IN3(n10625), .QN(
        \fadd_0_0_0_0_9/sub_784/B[1] ) );
  OAI21X1 U3170 ( .IN1(n10419), .IN2(n11597), .IN3(n11920), .QN(n10625) );
  NAND4X0 U3173 ( .IN1(n11919), .IN2(n11920), .IN3(n11921), .IN4(n11922), .QN(
        n10419) );
  AO22X1 U3174 ( .IN1(n14312), .IN2(n13513), .IN3(n10617), .IN4(n13626), .Q(
        \fadd_0_0_0_0_9/newy_11 ) );
  AO22X1 U3175 ( .IN1(n14312), .IN2(n13504), .IN3(n10617), .IN4(n13893), .Q(
        \fadd_0_0_0_0_9/newy_10 ) );
  AO22X1 U3176 ( .IN1(n14312), .IN2(n5338), .IN3(n10617), .IN4(n5350), .Q(
        \fadd_0_0_0_0_9/newx [8]) );
  AO22X1 U3179 ( .IN1(n14312), .IN2(n5337), .IN3(n10617), .IN4(n5349), .Q(
        \fadd_0_0_0_0_9/newx [7]) );
  AO22X1 U3182 ( .IN1(n14312), .IN2(n5336), .IN3(n10617), .IN4(n5348), .Q(
        \fadd_0_0_0_0_9/newx [6]) );
  AO22X1 U3185 ( .IN1(n14312), .IN2(n5335), .IN3(n10617), .IN4(n5347), .Q(
        \fadd_0_0_0_0_9/newx [5]) );
  AO22X1 U3188 ( .IN1(n14312), .IN2(n5334), .IN3(n10617), .IN4(n5346), .Q(
        \fadd_0_0_0_0_9/newx [4]) );
  AO22X1 U3191 ( .IN1(n14312), .IN2(n13712), .IN3(n10617), .IN4(n13574), .Q(
        \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ) );
  AO22X1 U3194 ( .IN1(n14312), .IN2(n13690), .IN3(n10617), .IN4(n13557), .Q(
        \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ) );
  AO22X1 U3197 ( .IN1(n14312), .IN2(n13669), .IN3(n10617), .IN4(n13532), .Q(
        \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ) );
  AO22X1 U3201 ( .IN1(n14312), .IN2(n13893), .IN3(n10617), .IN4(n13504), .Q(
        \fadd_0_0_0_0_9/newx [10]) );
  AO22X1 U3203 ( .IN1(n14312), .IN2(n13641), .IN3(n10617), .IN4(n13521), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ) );
  XOR2X1 U3206 ( .IN1(n10627), .IN2(n14879), .Q(
        \fadd_0_0_0_0_9/fracyfarxorop [6]) );
  XOR2X1 U3208 ( .IN1(n10630), .IN2(n12782), .Q(
        \fadd_0_0_0_0_9/fracyfarxorop [5]) );
  OA21X1 U3209 ( .IN1(n12779), .IN2(n14881), .IN3(n14876), .Q(n10630) );
  XOR2X1 U3211 ( .IN1(n10633), .IN2(n12782), .Q(
        \fadd_0_0_0_0_9/fracyfarxorop [4]) );
  OA22X1 U3212 ( .IN1(n14878), .IN2(n10634), .IN3(n12779), .IN4(n10635), .Q(
        n10633) );
  AO22X1 U3214 ( .IN1(n10637), .IN2(n14878), .IN3(n10638), .IN4(n12779), .Q(
        \fadd_0_0_0_0_9/fracyfarxorop [3]) );
  XOR2X1 U3215 ( .IN1(n10635), .IN2(n12782), .Q(n10638) );
  AO21X1 U3216 ( .IN1(n14882), .IN2(n10640), .IN3(n14875), .Q(n10635) );
  AO22X1 U3217 ( .IN1(n10642), .IN2(n14878), .IN3(n10637), .IN4(n12779), .Q(
        \fadd_0_0_0_0_9/fracyfarxorop [2]) );
  XOR2X1 U3218 ( .IN1(n14879), .IN2(n10643), .Q(n10637) );
  OA22X1 U3219 ( .IN1(n10636), .IN2(n10644), .IN3(n10645), .IN4(n10632), .Q(
        n10643) );
  AO22X1 U3221 ( .IN1(n10647), .IN2(n14878), .IN3(n10642), .IN4(n12779), .Q(
        \fadd_0_0_0_0_9/fracyfarxorop [1]) );
  XOR2X1 U3222 ( .IN1(n14879), .IN2(n10648), .Q(n10642) );
  OA22X1 U3223 ( .IN1(n10649), .IN2(n10644), .IN3(n14877), .IN4(n10650), .Q(
        n10648) );
  AO22X1 U3225 ( .IN1(n10647), .IN2(n12779), .IN3(n10651), .IN4(n14878), .Q(
        \fadd_0_0_0_0_9/fracyfarxorop [0]) );
  XOR2X1 U3227 ( .IN1(n12780), .IN2(n12782), .Q(n10651) );
  OA22X1 U3228 ( .IN1(n14877), .IN2(n12781), .IN3(n14884), .IN4(n14874), .Q(
        n12780) );
  XOR2X1 U3232 ( .IN1(n14879), .IN2(n10653), .Q(n10647) );
  AOI22X1 U3233 ( .IN1(n14883), .IN2(n14875), .IN3(n10646), .IN4(
        \fadd_0_0_0_0_9/rightshiftercomponent/level2[1] ), .QN(n10653) );
  OA221X1 U3237 ( .IN1(n14886), .IN2(n14312), .IN3(n14888), .IN4(n10617), 
        .IN5(n10652), .Q(n10640) );
  OA221X1 U3241 ( .IN1(n14887), .IN2(n14312), .IN3(n14889), .IN4(n10617), 
        .IN5(n10652), .Q(n10646) );
  OA22X1 U3242 ( .IN1(n14312), .IN2(n10616), .IN3(n10620), .IN4(n10617), .Q(
        n10652) );
  XOR2X1 U3248 ( .IN1(n14880), .IN2(\fadd_0_0_0_0_9/newy_9 ), .Q(n12782) );
  AO22X1 U3249 ( .IN1(n14312), .IN2(n13583), .IN3(n10617), .IN4(n13721), .Q(
        \fadd_0_0_0_0_9/newy_9 ) );
  OA22X1 U3253 ( .IN1(n10617), .IN2(n11833), .IN3(n14312), .IN4(n11844), .Q(
        n10611) );
  AO22X1 U3255 ( .IN1(n14885), .IN2(n14882), .IN3(n14881), .IN4(n10654), .Q(
        \fadd_0_0_0_0_9/fracyclose1 [3]) );
  OA22X1 U3257 ( .IN1(n10617), .IN2(n11838), .IN3(n14312), .IN4(n11827), .Q(
        n10636) );
  AO22X1 U3258 ( .IN1(n14885), .IN2(n14883), .IN3(n14882), .IN4(n10654), .Q(
        \fadd_0_0_0_0_9/fracyclose1 [2]) );
  OA22X1 U3260 ( .IN1(n10617), .IN2(n11837), .IN3(n14312), .IN4(n11826), .Q(
        n10649) );
  AO22X1 U3261 ( .IN1(n14883), .IN2(n10654), .IN3(n14885), .IN4(n14884), .Q(
        \fadd_0_0_0_0_9/fracyclose1 [1]) );
  OA22X1 U3264 ( .IN1(n10617), .IN2(n11836), .IN3(n14312), .IN4(n11825), .Q(
        n10645) );
  OA22X1 U3266 ( .IN1(n10617), .IN2(n11835), .IN3(n14312), .IN4(n11824), .Q(
        n10655) );
  AO22X1 U3268 ( .IN1(\fadd_0_0_0_0_9/exponentdifferenceyx [0]), .IN2(n14312), 
        .IN3(\fadd_0_0_0_0_9/exponentdifferencexy [0]), .IN4(n10617), .Q(
        n10654) );
  OA22X1 U3271 ( .IN1(n11834), .IN2(n10658), .IN3(
        \fadd_0_0_0_0_9/sub_707/carry [5]), .IN4(n13504), .Q(n10657) );
  AO22X1 U3278 ( .IN1(\fadd_0_0_0_0_9/fracrcloseymx [5]), .IN2(n14114), .IN3(
        \fadd_0_0_0_0_9/fracrclosexmy [5]), .IN4(n14649), .Q(
        \fadd_0_0_0_0_9/fracrclose1 [5]) );
  AO22X1 U3279 ( .IN1(\fadd_0_0_0_0_9/fracrcloseymx [4]), .IN2(n14114), .IN3(
        \fadd_0_0_0_0_9/fracrclosexmy [4]), .IN4(n14649), .Q(
        \fadd_0_0_0_0_9/fracrclose1 [4]) );
  AO22X1 U3280 ( .IN1(\fadd_0_0_0_0_9/fracrcloseymx [3]), .IN2(n14114), .IN3(
        \fadd_0_0_0_0_9/fracrclosexmy [3]), .IN4(n14649), .Q(
        \fadd_0_0_0_0_9/fracrclose1 [3]) );
  AO22X1 U3281 ( .IN1(\fadd_0_0_0_0_9/fracrcloseymx [2]), .IN2(n14114), .IN3(
        \fadd_0_0_0_0_9/fracrclosexmy [2]), .IN4(n14649), .Q(
        \fadd_0_0_0_0_9/fracrclose1 [2]) );
  AO22X1 U3282 ( .IN1(\fadd_0_0_0_0_9/fracrcloseymx [1]), .IN2(n14114), .IN3(
        \fadd_0_0_0_0_9/fracrclosexmy [1]), .IN4(n14649), .Q(
        \fadd_0_0_0_0_9/fracrclose1 [1]) );
  AO22X1 U3283 ( .IN1(\fadd_0_0_0_0_9/fracrcloseymx [0]), .IN2(n14114), .IN3(
        \fadd_0_0_0_0_9/fracrcloseymx [0]), .IN4(n14649), .Q(
        \fadd_0_0_0_0_9/fracrclose1 [0]) );
  NOR3X0 U3287 ( .IN1(n14960), .IN2(n11596), .IN3(n10593), .QN(
        \fadd_0_0_0_0_9/cinaddfar ) );
  AND2X1 U3288 ( .IN1(\fadd_0_0_0_0_9/rightshiftercomponent/level1_d2[0] ), 
        .IN2(\fadd_0_0_0_0_9/rightshiftercomponent/ps_d2[0] ), .Q(n10593) );
  NOR3X0 U3290 ( .IN1(n14936), .IN2(n11594), .IN3(n10418), .QN(
        \fadd_0_0_0_0_8/zerofromclose ) );
  NAND3X0 U3292 ( .IN1(n13671), .IN2(n13482), .IN3(n10667), .QN(n10664) );
  NAND3X0 U3293 ( .IN1(n10668), .IN2(n10669), .IN3(n12846), .QN(n10663) );
  AO222X1 U3298 ( .IN1(\fadd_0_0_0_0_8/fracresultfar0 [1]), .IN2(n14870), 
        .IN3(\fadd_0_0_0_0_8/fracresultfar0 [2]), .IN4(n10673), .IN5(
        \fadd_0_0_0_0_8/fracresultfar0 [0]), .IN6(
        \fadd_0_0_0_0_8/add_859/B[1] ), .Q(n10668) );
  AO22X1 U3299 ( .IN1(n10677), .IN2(
        \fadd_0_0_0_0_8/rightshiftercomponent/ps_d1 [1]), .IN3(n10678), .IN4(
        \fadd_0_0_0_0_8/rightshiftercomponent/ps_d1 [2]), .Q(
        \fadd_0_0_0_0_8/rightshiftercomponent/n389_o ) );
  AO22X1 U3302 ( .IN1(n13643), .IN2(\fadd_0_0_0_0_8/exponentresultclose_d1 [5]), .IN3(\fadd_0_0_0_0_8/exponentresultfar1 [5]), .IN4(n12846), .Q(
        \fadd_0_0_0_0_8/resultbeforeround [9]) );
  AO22X1 U3303 ( .IN1(n13643), .IN2(\fadd_0_0_0_0_8/exponentresultclose_d1 [4]), .IN3(\fadd_0_0_0_0_8/exponentresultfar1 [4]), .IN4(n12846), .Q(
        \fadd_0_0_0_0_8/resultbeforeround [8]) );
  AO22X1 U3304 ( .IN1(n13643), .IN2(\fadd_0_0_0_0_8/exponentresultclose_d1 [3]), .IN3(\fadd_0_0_0_0_8/exponentresultfar1 [3]), .IN4(n12846), .Q(
        \fadd_0_0_0_0_8/resultbeforeround [7]) );
  AO22X1 U3305 ( .IN1(n13643), .IN2(\fadd_0_0_0_0_8/exponentresultclose_d1 [2]), .IN3(\fadd_0_0_0_0_8/exponentresultfar1 [2]), .IN4(n12846), .Q(
        \fadd_0_0_0_0_8/resultbeforeround [6]) );
  AO22X1 U3306 ( .IN1(n13643), .IN2(\fadd_0_0_0_0_8/exponentresultclose_d1 [1]), .IN3(\fadd_0_0_0_0_8/exponentresultfar1 [1]), .IN4(n12846), .Q(
        \fadd_0_0_0_0_8/resultbeforeround [5]) );
  AO22X1 U3307 ( .IN1(n13643), .IN2(\fadd_0_0_0_0_8/exponentresultclose_d1 [0]), .IN3(\fadd_0_0_0_0_8/exponentresultfar1 [0]), .IN4(n12846), .Q(
        \fadd_0_0_0_0_8/resultbeforeround [4]) );
  AO222X1 U3308 ( .IN1(n10667), .IN2(\fadd_0_0_0_0_8/norm/level1_d1[4] ), 
        .IN3(n10680), .IN4(n13692), .IN5(n12846), .IN6(n10682), .Q(
        \fadd_0_0_0_0_8/resultbeforeround [3]) );
  AO222X1 U3309 ( .IN1(\fadd_0_0_0_0_8/fracresultfar0 [5]), .IN2(n14870), 
        .IN3(n10673), .IN4(\fadd_0_0_0_0_8/fracresultfar0 [6]), .IN5(
        \fadd_0_0_0_0_8/fracresultfar0 [4]), .IN6(
        \fadd_0_0_0_0_8/add_859/B[1] ), .Q(n10682) );
  AO222X1 U3310 ( .IN1(n10667), .IN2(n13692), .IN3(n10680), .IN4(n13550), 
        .IN5(n12846), .IN6(n10684), .Q(\fadd_0_0_0_0_8/resultbeforeround [2])
         );
  AO222X1 U3311 ( .IN1(\fadd_0_0_0_0_8/fracresultfar0 [4]), .IN2(n14870), 
        .IN3(\fadd_0_0_0_0_8/fracresultfar0 [5]), .IN4(n10673), .IN5(
        \fadd_0_0_0_0_8/add_859/B[1] ), .IN6(
        \fadd_0_0_0_0_8/fracresultfar0 [3]), .Q(n10684) );
  AO222X1 U3313 ( .IN1(n10667), .IN2(n13550), .IN3(n10680), .IN4(n13482), 
        .IN5(n12846), .IN6(n10685), .Q(\fadd_0_0_0_0_8/resultbeforeround [1])
         );
  AO222X1 U3314 ( .IN1(\fadd_0_0_0_0_8/fracresultfar0 [3]), .IN2(n14870), 
        .IN3(\fadd_0_0_0_0_8/fracresultfar0 [4]), .IN4(n10673), .IN5(
        \fadd_0_0_0_0_8/add_859/B[1] ), .IN6(
        \fadd_0_0_0_0_8/fracresultfar0 [2]), .Q(n10685) );
  AO22X1 U3316 ( .IN1(n13643), .IN2(\fadd_0_0_0_0_8/exponentresultclose_d1 [6]), .IN3(\fadd_0_0_0_0_8/exponentresultfar1 [6]), .IN4(n12846), .Q(
        \fadd_0_0_0_0_8/resultbeforeround [10]) );
  AO222X1 U3317 ( .IN1(n10667), .IN2(n13482), .IN3(n10680), .IN4(n13671), 
        .IN5(n12846), .IN6(n10675), .Q(\fadd_0_0_0_0_8/resultbeforeround [0])
         );
  AO222X1 U3318 ( .IN1(\fadd_0_0_0_0_8/fracresultfar0 [2]), .IN2(n14870), 
        .IN3(\fadd_0_0_0_0_8/fracresultfar0 [3]), .IN4(n10673), .IN5(
        \fadd_0_0_0_0_8/fracresultfar0 [1]), .IN6(
        \fadd_0_0_0_0_8/add_859/B[1] ), .Q(n10675) );
  AND2X1 U3325 ( .IN1(n12865), .IN2(n13643), .Q(n10667) );
  OA221X1 U3327 ( .IN1(n10686), .IN2(n10687), .IN3(n10688), .IN4(n10689), 
        .IN5(n10690), .Q(\fadd_0_0_0_0_8/ressign ) );
  XOR2X1 U3328 ( .IN1(n10691), .IN2(n10692), .Q(n10690) );
  OR3X1 U3329 ( .IN1(\fadd_0_0_0_0_8/fracrcloseymx [0]), .IN2(
        \fadd_0_0_0_0_8/fracrcloseymx [1]), .IN3(n10691), .Q(n10689) );
  OR4X1 U3332 ( .IN1(\fadd_0_0_0_0_8/fracrcloseymx [2]), .IN2(
        \fadd_0_0_0_0_8/fracrcloseymx [3]), .IN3(
        \fadd_0_0_0_0_8/fracrcloseymx [4]), .IN4(
        \fadd_0_0_0_0_8/fracrcloseymx [5]), .Q(n10688) );
  OR4X1 U3333 ( .IN1(n10693), .IN2(\fadd_0_0_0_0_8/fracrcloseymx [0]), .IN3(
        \fadd_0_0_0_0_8/fracrclosexmy [1]), .IN4(
        \fadd_0_0_0_0_8/fracrclosexmy [2]), .Q(n10687) );
  AO21X1 U3334 ( .IN1(n10694), .IN2(n10695), .IN3(n14847), .Q(n10693) );
  NAND4X0 U3335 ( .IN1(n10697), .IN2(n10698), .IN3(n14855), .IN4(n14854), .QN(
        n10695) );
  NAND4X0 U3336 ( .IN1(n10701), .IN2(n14311), .IN3(n14857), .IN4(n14856), .QN(
        n10694) );
  AO21X1 U3338 ( .IN1(\fadd_0_0_0_0_8/sub_784/B[1] ), .IN2(n14056), .IN3(
        n10706), .Q(\fadd_0_0_0_0_8/norm/level1 [4]) );
  OAI22X1 U3340 ( .IN1(n14936), .IN2(n11585), .IN3(n10707), .IN4(n11917), .QN(
        \fadd_0_0_0_0_8/norm/level1 [3]) );
  OAI22X1 U3341 ( .IN1(n14936), .IN2(n11584), .IN3(n10707), .IN4(n11918), .QN(
        \fadd_0_0_0_0_8/norm/level1 [2]) );
  NOR3X0 U3346 ( .IN1(n13540), .IN2(n8664), .IN3(n10706), .QN(
        \fadd_0_0_0_0_8/sub_784/B[1] ) );
  OAI21X1 U3347 ( .IN1(n10418), .IN2(n11584), .IN3(n11916), .QN(n10706) );
  NAND4X0 U3350 ( .IN1(n11915), .IN2(n11916), .IN3(n11917), .IN4(n11918), .QN(
        n10418) );
  AO22X1 U3351 ( .IN1(n14311), .IN2(n13630), .IN3(n10698), .IN4(n13501), .Q(
        \fadd_0_0_0_0_8/newy_11 ) );
  AO22X1 U3352 ( .IN1(n14311), .IN2(n13628), .IN3(n10698), .IN4(n13588), .Q(
        \fadd_0_0_0_0_8/newy_10 ) );
  OAI22X1 U3353 ( .IN1(n10698), .IN2(n14619), .IN3(n14311), .IN4(n14624), .QN(
        \fadd_0_0_0_0_8/newx [8]) );
  OAI22X1 U3354 ( .IN1(n10698), .IN2(n14620), .IN3(n14311), .IN4(n14625), .QN(
        \fadd_0_0_0_0_8/newx [7]) );
  OAI22X1 U3355 ( .IN1(n10698), .IN2(n14621), .IN3(n14311), .IN4(n14626), .QN(
        \fadd_0_0_0_0_8/newx [6]) );
  OAI22X1 U3356 ( .IN1(n10698), .IN2(n14622), .IN3(n14311), .IN4(n14627), .QN(
        \fadd_0_0_0_0_8/newx [5]) );
  OAI22X1 U3357 ( .IN1(n10698), .IN2(n14623), .IN3(n14311), .IN4(n14628), .QN(
        \fadd_0_0_0_0_8/newx [4]) );
  OAI22X1 U3359 ( .IN1(n10698), .IN2(n11858), .IN3(n14311), .IN4(n11870), .QN(
        \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ) );
  AO22X1 U3362 ( .IN1(n14311), .IN2(n13588), .IN3(n10698), .IN4(n13628), .Q(
        \fadd_0_0_0_0_8/newx [10]) );
  OAI22X1 U3364 ( .IN1(n10698), .IN2(n11856), .IN3(n14311), .IN4(n11868), .QN(
        \add_0_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ) );
  XOR2X1 U3365 ( .IN1(n10710), .IN2(n14847), .Q(
        \fadd_0_0_0_0_8/fracyfarxorop [6]) );
  XOR2X1 U3367 ( .IN1(n10713), .IN2(n12772), .Q(
        \fadd_0_0_0_0_8/fracyfarxorop [5]) );
  OA21X1 U3368 ( .IN1(n12769), .IN2(n14849), .IN3(n14844), .Q(n10713) );
  XOR2X1 U3370 ( .IN1(n10716), .IN2(n12772), .Q(
        \fadd_0_0_0_0_8/fracyfarxorop [4]) );
  OA22X1 U3371 ( .IN1(n14846), .IN2(n10717), .IN3(n12769), .IN4(n10718), .Q(
        n10716) );
  AO22X1 U3373 ( .IN1(n10720), .IN2(n14846), .IN3(n10721), .IN4(n12769), .Q(
        \fadd_0_0_0_0_8/fracyfarxorop [3]) );
  XOR2X1 U3374 ( .IN1(n10718), .IN2(n12772), .Q(n10721) );
  AO21X1 U3375 ( .IN1(n14850), .IN2(n10723), .IN3(n14843), .Q(n10718) );
  AO22X1 U3376 ( .IN1(n10725), .IN2(n14846), .IN3(n10720), .IN4(n12769), .Q(
        \fadd_0_0_0_0_8/fracyfarxorop [2]) );
  XOR2X1 U3377 ( .IN1(n14847), .IN2(n10726), .Q(n10720) );
  OA22X1 U3378 ( .IN1(n10719), .IN2(n10727), .IN3(n10728), .IN4(n10715), .Q(
        n10726) );
  AO22X1 U3380 ( .IN1(n10730), .IN2(n14846), .IN3(n10725), .IN4(n12769), .Q(
        \fadd_0_0_0_0_8/fracyfarxorop [1]) );
  XOR2X1 U3381 ( .IN1(n14847), .IN2(n10731), .Q(n10725) );
  OA22X1 U3382 ( .IN1(n10732), .IN2(n10727), .IN3(n14845), .IN4(n10733), .Q(
        n10731) );
  AO22X1 U3384 ( .IN1(n10730), .IN2(n12769), .IN3(n10734), .IN4(n14846), .Q(
        \fadd_0_0_0_0_8/fracyfarxorop [0]) );
  XOR2X1 U3386 ( .IN1(n12770), .IN2(n12772), .Q(n10734) );
  OA22X1 U3387 ( .IN1(n14845), .IN2(n12771), .IN3(n14852), .IN4(n14842), .Q(
        n12770) );
  XOR2X1 U3391 ( .IN1(n14847), .IN2(n10736), .Q(n10730) );
  AOI22X1 U3392 ( .IN1(n14851), .IN2(n14843), .IN3(n10729), .IN4(
        \fadd_0_0_0_0_8/rightshiftercomponent/level2[1] ), .QN(n10736) );
  OA221X1 U3396 ( .IN1(n14854), .IN2(n14311), .IN3(n14856), .IN4(n10698), 
        .IN5(n10735), .Q(n10723) );
  OA221X1 U3400 ( .IN1(n14855), .IN2(n14311), .IN3(n14857), .IN4(n10698), 
        .IN5(n10735), .Q(n10729) );
  OA22X1 U3401 ( .IN1(n14311), .IN2(n10697), .IN3(n10701), .IN4(n10698), .Q(
        n10735) );
  XOR2X1 U3407 ( .IN1(n14848), .IN2(\fadd_0_0_0_0_8/newy_9 ), .Q(n12772) );
  OAI22X1 U3408 ( .IN1(n10698), .IN2(n11877), .IN3(n14311), .IN4(n11865), .QN(
        \fadd_0_0_0_0_8/newy_9 ) );
  OA22X1 U3410 ( .IN1(n10698), .IN2(n11865), .IN3(n14311), .IN4(n11877), .Q(
        n10692) );
  AO22X1 U3412 ( .IN1(n14853), .IN2(n14850), .IN3(n14849), .IN4(n10737), .Q(
        \fadd_0_0_0_0_8/fracyclose1 [3]) );
  OA22X1 U3414 ( .IN1(n10698), .IN2(n11871), .IN3(n14311), .IN4(n11859), .Q(
        n10719) );
  AO22X1 U3415 ( .IN1(n14853), .IN2(n14851), .IN3(n14850), .IN4(n10737), .Q(
        \fadd_0_0_0_0_8/fracyclose1 [2]) );
  OA22X1 U3417 ( .IN1(n10698), .IN2(n11870), .IN3(n14311), .IN4(n11858), .Q(
        n10732) );
  AO22X1 U3418 ( .IN1(n14851), .IN2(n10737), .IN3(n14853), .IN4(n14852), .Q(
        \fadd_0_0_0_0_8/fracyclose1 [1]) );
  OA22X1 U3421 ( .IN1(n10698), .IN2(n11869), .IN3(n14311), .IN4(n11857), .Q(
        n10728) );
  OA22X1 U3423 ( .IN1(n10698), .IN2(n11868), .IN3(n14311), .IN4(n11856), .Q(
        n10738) );
  AO22X1 U3425 ( .IN1(\fadd_0_0_0_0_8/exponentdifferenceyx [0]), .IN2(n14311), 
        .IN3(\fadd_0_0_0_0_8/exponentdifferencexy [0]), .IN4(n10698), .Q(
        n10737) );
  OA22X1 U3428 ( .IN1(n11867), .IN2(n10741), .IN3(
        \fadd_0_0_0_0_8/sub_707/carry [5]), .IN4(n13628), .Q(n10740) );
  AO22X1 U3435 ( .IN1(\fadd_0_0_0_0_8/fracrcloseymx [5]), .IN2(n14118), .IN3(
        \fadd_0_0_0_0_8/fracrclosexmy [5]), .IN4(n14650), .Q(
        \fadd_0_0_0_0_8/fracrclose1 [5]) );
  AO22X1 U3436 ( .IN1(\fadd_0_0_0_0_8/fracrcloseymx [4]), .IN2(n14118), .IN3(
        \fadd_0_0_0_0_8/fracrclosexmy [4]), .IN4(n14650), .Q(
        \fadd_0_0_0_0_8/fracrclose1 [4]) );
  AO22X1 U3437 ( .IN1(\fadd_0_0_0_0_8/fracrcloseymx [3]), .IN2(n14118), .IN3(
        \fadd_0_0_0_0_8/fracrclosexmy [3]), .IN4(n14650), .Q(
        \fadd_0_0_0_0_8/fracrclose1 [3]) );
  AO22X1 U3438 ( .IN1(\fadd_0_0_0_0_8/fracrcloseymx [2]), .IN2(n14118), .IN3(
        \fadd_0_0_0_0_8/fracrclosexmy [2]), .IN4(n14650), .Q(
        \fadd_0_0_0_0_8/fracrclose1 [2]) );
  AO22X1 U3439 ( .IN1(\fadd_0_0_0_0_8/fracrcloseymx [1]), .IN2(n14118), .IN3(
        \fadd_0_0_0_0_8/fracrclosexmy [1]), .IN4(n14650), .Q(
        \fadd_0_0_0_0_8/fracrclose1 [1]) );
  AO22X1 U3440 ( .IN1(\fadd_0_0_0_0_8/fracrcloseymx [0]), .IN2(n14118), .IN3(
        \fadd_0_0_0_0_8/fracrcloseymx [0]), .IN4(n14650), .Q(
        \fadd_0_0_0_0_8/fracrclose1 [0]) );
  NOR3X0 U3444 ( .IN1(n15002), .IN2(n11583), .IN3(n10674), .QN(
        \fadd_0_0_0_0_8/cinaddfar ) );
  AND2X1 U3445 ( .IN1(\fadd_0_0_0_0_8/rightshiftercomponent/level1_d2[0] ), 
        .IN2(\fadd_0_0_0_0_8/rightshiftercomponent/ps_d2[0] ), .Q(n10674) );
  NOR3X0 U3447 ( .IN1(n14935), .IN2(n11581), .IN3(n10417), .QN(
        \fadd_0_0_0_0_7/zerofromclose ) );
  NAND3X0 U3449 ( .IN1(n13683), .IN2(n13491), .IN3(n10750), .QN(n10747) );
  NAND3X0 U3450 ( .IN1(n10751), .IN2(n10752), .IN3(n12845), .QN(n10746) );
  AO222X1 U3455 ( .IN1(\fadd_0_0_0_0_7/fracresultfar0 [1]), .IN2(n14838), 
        .IN3(\fadd_0_0_0_0_7/fracresultfar0 [2]), .IN4(n10756), .IN5(
        \fadd_0_0_0_0_7/fracresultfar0 [0]), .IN6(n14231), .Q(n10751) );
  AO22X1 U3456 ( .IN1(n10760), .IN2(
        \fadd_0_0_0_0_7/rightshiftercomponent/ps_d1 [1]), .IN3(n10761), .IN4(
        \fadd_0_0_0_0_7/rightshiftercomponent/ps_d1 [2]), .Q(
        \fadd_0_0_0_0_7/rightshiftercomponent/n389_o ) );
  AO22X1 U3459 ( .IN1(n13652), .IN2(\fadd_0_0_0_0_7/exponentresultclose_d1 [5]), .IN3(\fadd_0_0_0_0_7/exponentresultfar1 [5]), .IN4(n12845), .Q(
        \fadd_0_0_0_0_7/resultbeforeround [9]) );
  AO22X1 U3460 ( .IN1(n13652), .IN2(\fadd_0_0_0_0_7/exponentresultclose_d1 [4]), .IN3(\fadd_0_0_0_0_7/exponentresultfar1 [4]), .IN4(n12845), .Q(
        \fadd_0_0_0_0_7/resultbeforeround [8]) );
  AO22X1 U3461 ( .IN1(n13652), .IN2(\fadd_0_0_0_0_7/exponentresultclose_d1 [3]), .IN3(\fadd_0_0_0_0_7/exponentresultfar1 [3]), .IN4(n12845), .Q(
        \fadd_0_0_0_0_7/resultbeforeround [7]) );
  AO22X1 U3462 ( .IN1(n13652), .IN2(\fadd_0_0_0_0_7/exponentresultclose_d1 [2]), .IN3(\fadd_0_0_0_0_7/exponentresultfar1 [2]), .IN4(n12845), .Q(
        \fadd_0_0_0_0_7/resultbeforeround [6]) );
  AO22X1 U3463 ( .IN1(n13652), .IN2(\fadd_0_0_0_0_7/exponentresultclose_d1 [1]), .IN3(\fadd_0_0_0_0_7/exponentresultfar1 [1]), .IN4(n12845), .Q(
        \fadd_0_0_0_0_7/resultbeforeround [5]) );
  AO22X1 U3464 ( .IN1(n13652), .IN2(\fadd_0_0_0_0_7/exponentresultclose_d1 [0]), .IN3(\fadd_0_0_0_0_7/exponentresultfar1 [0]), .IN4(n12845), .Q(
        \fadd_0_0_0_0_7/resultbeforeround [4]) );
  AO222X1 U3465 ( .IN1(n10750), .IN2(\fadd_0_0_0_0_7/norm/level1_d1[4] ), 
        .IN3(n10763), .IN4(n13704), .IN5(n12845), .IN6(n10765), .Q(
        \fadd_0_0_0_0_7/resultbeforeround [3]) );
  AO222X1 U3466 ( .IN1(\fadd_0_0_0_0_7/fracresultfar0 [5]), .IN2(n14838), 
        .IN3(n10756), .IN4(\fadd_0_0_0_0_7/fracresultfar0 [6]), .IN5(
        \fadd_0_0_0_0_7/fracresultfar0 [4]), .IN6(n14231), .Q(n10765) );
  AO222X1 U3467 ( .IN1(n10750), .IN2(n13704), .IN3(n10763), .IN4(n13568), 
        .IN5(n12845), .IN6(n10767), .Q(\fadd_0_0_0_0_7/resultbeforeround [2])
         );
  AO222X1 U3468 ( .IN1(\fadd_0_0_0_0_7/fracresultfar0 [4]), .IN2(n14838), 
        .IN3(\fadd_0_0_0_0_7/fracresultfar0 [5]), .IN4(n10756), .IN5(n14231), 
        .IN6(\fadd_0_0_0_0_7/fracresultfar0 [3]), .Q(n10767) );
  AO222X1 U3470 ( .IN1(n10750), .IN2(n13568), .IN3(n10763), .IN4(n13491), 
        .IN5(n12845), .IN6(n10768), .Q(\fadd_0_0_0_0_7/resultbeforeround [1])
         );
  AO222X1 U3471 ( .IN1(\fadd_0_0_0_0_7/fracresultfar0 [3]), .IN2(n14838), 
        .IN3(\fadd_0_0_0_0_7/fracresultfar0 [4]), .IN4(n10756), .IN5(n14231), 
        .IN6(\fadd_0_0_0_0_7/fracresultfar0 [2]), .Q(n10768) );
  AO22X1 U3473 ( .IN1(n13652), .IN2(\fadd_0_0_0_0_7/exponentresultclose_d1 [6]), .IN3(\fadd_0_0_0_0_7/exponentresultfar1 [6]), .IN4(n12845), .Q(
        \fadd_0_0_0_0_7/resultbeforeround [10]) );
  AO222X1 U3474 ( .IN1(n10750), .IN2(n13491), .IN3(n10763), .IN4(n13683), 
        .IN5(n12845), .IN6(n10758), .Q(\fadd_0_0_0_0_7/resultbeforeround [0])
         );
  AO222X1 U3475 ( .IN1(\fadd_0_0_0_0_7/fracresultfar0 [2]), .IN2(n14838), 
        .IN3(\fadd_0_0_0_0_7/fracresultfar0 [3]), .IN4(n10756), .IN5(
        \fadd_0_0_0_0_7/fracresultfar0 [1]), .IN6(n14231), .Q(n10758) );
  AND2X1 U3482 ( .IN1(n12863), .IN2(n13652), .Q(n10750) );
  OA221X1 U3484 ( .IN1(n10769), .IN2(n10770), .IN3(n10771), .IN4(n10772), 
        .IN5(n10773), .Q(\fadd_0_0_0_0_7/ressign ) );
  XOR2X1 U3485 ( .IN1(n10774), .IN2(n10775), .Q(n10773) );
  OR3X1 U3486 ( .IN1(\fadd_0_0_0_0_7/fracrcloseymx [0]), .IN2(
        \fadd_0_0_0_0_7/fracrcloseymx [1]), .IN3(n10774), .Q(n10772) );
  OR4X1 U3489 ( .IN1(\fadd_0_0_0_0_7/fracrcloseymx [2]), .IN2(
        \fadd_0_0_0_0_7/fracrcloseymx [3]), .IN3(
        \fadd_0_0_0_0_7/fracrcloseymx [4]), .IN4(
        \fadd_0_0_0_0_7/fracrcloseymx [5]), .Q(n10771) );
  OR4X1 U3490 ( .IN1(n10776), .IN2(\fadd_0_0_0_0_7/fracrcloseymx [0]), .IN3(
        \fadd_0_0_0_0_7/fracrclosexmy [1]), .IN4(
        \fadd_0_0_0_0_7/fracrclosexmy [2]), .Q(n10770) );
  AO21X1 U3491 ( .IN1(n10777), .IN2(n10778), .IN3(n14826), .Q(n10776) );
  NAND4X0 U3492 ( .IN1(n10780), .IN2(n10781), .IN3(n14834), .IN4(n14833), .QN(
        n10778) );
  NAND4X0 U3493 ( .IN1(n10784), .IN2(n14310), .IN3(n14836), .IN4(n14835), .QN(
        n10777) );
  AO21X1 U3495 ( .IN1(\fadd_0_0_0_0_7/sub_784/B[1] ), .IN2(n14055), .IN3(
        n10789), .Q(\fadd_0_0_0_0_7/norm/level1 [4]) );
  OAI22X1 U3497 ( .IN1(n14935), .IN2(n11572), .IN3(n10790), .IN4(n11913), .QN(
        \fadd_0_0_0_0_7/norm/level1 [3]) );
  OAI22X1 U3498 ( .IN1(n14935), .IN2(n11571), .IN3(n10790), .IN4(n11914), .QN(
        \fadd_0_0_0_0_7/norm/level1 [2]) );
  NOR3X0 U3503 ( .IN1(n13541), .IN2(n8660), .IN3(n10789), .QN(
        \fadd_0_0_0_0_7/sub_784/B[1] ) );
  OAI21X1 U3504 ( .IN1(n10417), .IN2(n11571), .IN3(n11912), .QN(n10789) );
  NAND4X0 U3507 ( .IN1(n11911), .IN2(n11912), .IN3(n11913), .IN4(n11914), .QN(
        n10417) );
  AO22X1 U3508 ( .IN1(n14310), .IN2(n13512), .IN3(n10781), .IN4(n13625), .Q(
        \fadd_0_0_0_0_7/newy_11 ) );
  AO22X1 U3509 ( .IN1(n14310), .IN2(n13475), .IN3(n10781), .IN4(n13892), .Q(
        \fadd_0_0_0_0_7/newy_10 ) );
  AO22X1 U3510 ( .IN1(n14310), .IN2(n5482), .IN3(n10781), .IN4(n5494), .Q(
        \fadd_0_0_0_0_7/newx [8]) );
  AO22X1 U3513 ( .IN1(n14310), .IN2(n5481), .IN3(n10781), .IN4(n5493), .Q(
        \fadd_0_0_0_0_7/newx [7]) );
  AO22X1 U3516 ( .IN1(n14310), .IN2(n5480), .IN3(n10781), .IN4(n5492), .Q(
        \fadd_0_0_0_0_7/newx [6]) );
  AO22X1 U3519 ( .IN1(n14310), .IN2(n5479), .IN3(n10781), .IN4(n5491), .Q(
        \fadd_0_0_0_0_7/newx [5]) );
  AO22X1 U3522 ( .IN1(n14310), .IN2(n5478), .IN3(n10781), .IN4(n5490), .Q(
        \fadd_0_0_0_0_7/newx [4]) );
  AO22X1 U3525 ( .IN1(n14310), .IN2(n13711), .IN3(n10781), .IN4(n13573), .Q(
        \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ) );
  AO22X1 U3528 ( .IN1(n14310), .IN2(n13689), .IN3(n10781), .IN4(n13556), .Q(
        \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ) );
  AO22X1 U3531 ( .IN1(n14310), .IN2(n13668), .IN3(n10781), .IN4(n13531), .Q(
        \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ) );
  AO22X1 U3535 ( .IN1(n14310), .IN2(n13892), .IN3(n10781), .IN4(n13475), .Q(
        \fadd_0_0_0_0_7/newx [10]) );
  AO22X1 U3537 ( .IN1(n14310), .IN2(n13640), .IN3(n10781), .IN4(n13520), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ) );
  XOR2X1 U3540 ( .IN1(n10791), .IN2(n14826), .Q(
        \fadd_0_0_0_0_7/fracyfarxorop [6]) );
  XOR2X1 U3542 ( .IN1(n10794), .IN2(n12762), .Q(
        \fadd_0_0_0_0_7/fracyfarxorop [5]) );
  OA21X1 U3543 ( .IN1(n12759), .IN2(n14828), .IN3(n14823), .Q(n10794) );
  XOR2X1 U3545 ( .IN1(n10797), .IN2(n12762), .Q(
        \fadd_0_0_0_0_7/fracyfarxorop [4]) );
  OA22X1 U3546 ( .IN1(n14825), .IN2(n10798), .IN3(n12759), .IN4(n10799), .Q(
        n10797) );
  AO22X1 U3548 ( .IN1(n10801), .IN2(n14825), .IN3(n10802), .IN4(n12759), .Q(
        \fadd_0_0_0_0_7/fracyfarxorop [3]) );
  XOR2X1 U3549 ( .IN1(n10799), .IN2(n12762), .Q(n10802) );
  AO21X1 U3550 ( .IN1(n14829), .IN2(n10804), .IN3(n14822), .Q(n10799) );
  AO22X1 U3551 ( .IN1(n10806), .IN2(n14825), .IN3(n10801), .IN4(n12759), .Q(
        \fadd_0_0_0_0_7/fracyfarxorop [2]) );
  XOR2X1 U3552 ( .IN1(n14826), .IN2(n10807), .Q(n10801) );
  OA22X1 U3553 ( .IN1(n10800), .IN2(n10808), .IN3(n10809), .IN4(n10796), .Q(
        n10807) );
  AO22X1 U3555 ( .IN1(n10811), .IN2(n14825), .IN3(n10806), .IN4(n12759), .Q(
        \fadd_0_0_0_0_7/fracyfarxorop [1]) );
  XOR2X1 U3556 ( .IN1(n14826), .IN2(n10812), .Q(n10806) );
  OA22X1 U3557 ( .IN1(n10813), .IN2(n10808), .IN3(n14824), .IN4(n10814), .Q(
        n10812) );
  AO22X1 U3559 ( .IN1(n10811), .IN2(n12759), .IN3(n10815), .IN4(n14825), .Q(
        \fadd_0_0_0_0_7/fracyfarxorop [0]) );
  XOR2X1 U3561 ( .IN1(n12760), .IN2(n12762), .Q(n10815) );
  OA22X1 U3562 ( .IN1(n14824), .IN2(n12761), .IN3(n14831), .IN4(n14821), .Q(
        n12760) );
  XOR2X1 U3566 ( .IN1(n14826), .IN2(n10817), .Q(n10811) );
  AOI22X1 U3567 ( .IN1(n14830), .IN2(n14822), .IN3(n10810), .IN4(
        \fadd_0_0_0_0_7/rightshiftercomponent/level2[1] ), .QN(n10817) );
  OA221X1 U3571 ( .IN1(n14833), .IN2(n14310), .IN3(n14835), .IN4(n10781), 
        .IN5(n10816), .Q(n10804) );
  OA221X1 U3575 ( .IN1(n14834), .IN2(n14310), .IN3(n14836), .IN4(n10781), 
        .IN5(n10816), .Q(n10810) );
  OA22X1 U3576 ( .IN1(n14310), .IN2(n10780), .IN3(n10784), .IN4(n10781), .Q(
        n10816) );
  XOR2X1 U3582 ( .IN1(n14827), .IN2(\fadd_0_0_0_0_7/newy_9 ), .Q(n12762) );
  AO22X1 U3583 ( .IN1(n14310), .IN2(n13582), .IN3(n10781), .IN4(n13720), .Q(
        \fadd_0_0_0_0_7/newy_9 ) );
  OA22X1 U3587 ( .IN1(n10781), .IN2(n11749), .IN3(n14310), .IN4(n11760), .Q(
        n10775) );
  AO22X1 U3589 ( .IN1(n14832), .IN2(n14829), .IN3(n14828), .IN4(n10818), .Q(
        \fadd_0_0_0_0_7/fracyclose1 [3]) );
  OA22X1 U3591 ( .IN1(n10781), .IN2(n11754), .IN3(n14310), .IN4(n11743), .Q(
        n10800) );
  AO22X1 U3592 ( .IN1(n14832), .IN2(n14830), .IN3(n14829), .IN4(n10818), .Q(
        \fadd_0_0_0_0_7/fracyclose1 [2]) );
  OA22X1 U3594 ( .IN1(n10781), .IN2(n11753), .IN3(n14310), .IN4(n11742), .Q(
        n10813) );
  AO22X1 U3595 ( .IN1(n14830), .IN2(n10818), .IN3(n14832), .IN4(n14831), .Q(
        \fadd_0_0_0_0_7/fracyclose1 [1]) );
  OA22X1 U3598 ( .IN1(n10781), .IN2(n11752), .IN3(n14310), .IN4(n11741), .Q(
        n10809) );
  OA22X1 U3600 ( .IN1(n10781), .IN2(n11751), .IN3(n14310), .IN4(n11740), .Q(
        n10819) );
  AO22X1 U3602 ( .IN1(\fadd_0_0_0_0_7/exponentdifferenceyx [0]), .IN2(n14310), 
        .IN3(\fadd_0_0_0_0_7/exponentdifferencexy [0]), .IN4(n10781), .Q(
        n10818) );
  OA22X1 U3605 ( .IN1(n11750), .IN2(n10822), .IN3(
        \fadd_0_0_0_0_7/sub_707/carry [5]), .IN4(n13475), .Q(n10821) );
  AO22X1 U3612 ( .IN1(\fadd_0_0_0_0_7/fracrcloseymx [5]), .IN2(n14116), .IN3(
        \fadd_0_0_0_0_7/fracrclosexmy [5]), .IN4(n14645), .Q(
        \fadd_0_0_0_0_7/fracrclose1 [5]) );
  AO22X1 U3613 ( .IN1(\fadd_0_0_0_0_7/fracrcloseymx [4]), .IN2(n14116), .IN3(
        \fadd_0_0_0_0_7/fracrclosexmy [4]), .IN4(n14645), .Q(
        \fadd_0_0_0_0_7/fracrclose1 [4]) );
  AO22X1 U3614 ( .IN1(\fadd_0_0_0_0_7/fracrcloseymx [3]), .IN2(n14116), .IN3(
        \fadd_0_0_0_0_7/fracrclosexmy [3]), .IN4(n14645), .Q(
        \fadd_0_0_0_0_7/fracrclose1 [3]) );
  AO22X1 U3615 ( .IN1(\fadd_0_0_0_0_7/fracrcloseymx [2]), .IN2(n14116), .IN3(
        \fadd_0_0_0_0_7/fracrclosexmy [2]), .IN4(n14645), .Q(
        \fadd_0_0_0_0_7/fracrclose1 [2]) );
  AO22X1 U3616 ( .IN1(\fadd_0_0_0_0_7/fracrcloseymx [1]), .IN2(n14116), .IN3(
        \fadd_0_0_0_0_7/fracrclosexmy [1]), .IN4(n14645), .Q(
        \fadd_0_0_0_0_7/fracrclose1 [1]) );
  AO22X1 U3617 ( .IN1(\fadd_0_0_0_0_7/fracrcloseymx [0]), .IN2(n14116), .IN3(
        \fadd_0_0_0_0_7/fracrcloseymx [0]), .IN4(n14645), .Q(
        \fadd_0_0_0_0_7/fracrclose1 [0]) );
  NOR3X0 U3621 ( .IN1(n14951), .IN2(n11570), .IN3(n10757), .QN(
        \fadd_0_0_0_0_7/cinaddfar ) );
  AND2X1 U3622 ( .IN1(\fadd_0_0_0_0_7/rightshiftercomponent/level1_d2[0] ), 
        .IN2(\fadd_0_0_0_0_7/rightshiftercomponent/ps_d2[0] ), .Q(n10757) );
  NOR3X0 U3624 ( .IN1(n14934), .IN2(n11568), .IN3(n10416), .QN(
        \fadd_0_0_0_0_6/zerofromclose ) );
  NAND3X0 U3626 ( .IN1(n13678), .IN2(n13486), .IN3(n10831), .QN(n10828) );
  NAND3X0 U3627 ( .IN1(n10832), .IN2(n10833), .IN3(n12844), .QN(n10827) );
  AO222X1 U3632 ( .IN1(\fadd_0_0_0_0_6/fracresultfar0 [1]), .IN2(n14817), 
        .IN3(\fadd_0_0_0_0_6/fracresultfar0 [2]), .IN4(n10837), .IN5(
        \fadd_0_0_0_0_6/fracresultfar0 [0]), .IN6(
        \fadd_0_0_0_0_6/add_859/B[1] ), .Q(n10832) );
  AO22X1 U3633 ( .IN1(n10841), .IN2(
        \fadd_0_0_0_0_6/rightshiftercomponent/ps_d1 [1]), .IN3(n10842), .IN4(
        \fadd_0_0_0_0_6/rightshiftercomponent/ps_d1 [2]), .Q(
        \fadd_0_0_0_0_6/rightshiftercomponent/n389_o ) );
  AO22X1 U3636 ( .IN1(n13647), .IN2(\fadd_0_0_0_0_6/exponentresultclose_d1 [5]), .IN3(\fadd_0_0_0_0_6/exponentresultfar1 [5]), .IN4(n12844), .Q(
        \fadd_0_0_0_0_6/resultbeforeround [9]) );
  AO22X1 U3637 ( .IN1(n13647), .IN2(\fadd_0_0_0_0_6/exponentresultclose_d1 [4]), .IN3(\fadd_0_0_0_0_6/exponentresultfar1 [4]), .IN4(n12844), .Q(
        \fadd_0_0_0_0_6/resultbeforeround [8]) );
  AO22X1 U3638 ( .IN1(n13647), .IN2(\fadd_0_0_0_0_6/exponentresultclose_d1 [3]), .IN3(\fadd_0_0_0_0_6/exponentresultfar1 [3]), .IN4(n12844), .Q(
        \fadd_0_0_0_0_6/resultbeforeround [7]) );
  AO22X1 U3639 ( .IN1(n13647), .IN2(\fadd_0_0_0_0_6/exponentresultclose_d1 [2]), .IN3(\fadd_0_0_0_0_6/exponentresultfar1 [2]), .IN4(n12844), .Q(
        \fadd_0_0_0_0_6/resultbeforeround [6]) );
  AO22X1 U3640 ( .IN1(n13647), .IN2(\fadd_0_0_0_0_6/exponentresultclose_d1 [1]), .IN3(\fadd_0_0_0_0_6/exponentresultfar1 [1]), .IN4(n12844), .Q(
        \fadd_0_0_0_0_6/resultbeforeround [5]) );
  AO22X1 U3641 ( .IN1(n13647), .IN2(\fadd_0_0_0_0_6/exponentresultclose_d1 [0]), .IN3(\fadd_0_0_0_0_6/exponentresultfar1 [0]), .IN4(n12844), .Q(
        \fadd_0_0_0_0_6/resultbeforeround [4]) );
  AO222X1 U3642 ( .IN1(n10831), .IN2(\fadd_0_0_0_0_6/norm/level1_d1[4] ), 
        .IN3(n10844), .IN4(n13699), .IN5(n12844), .IN6(n10846), .Q(
        \fadd_0_0_0_0_6/resultbeforeround [3]) );
  AO222X1 U3643 ( .IN1(\fadd_0_0_0_0_6/fracresultfar0 [5]), .IN2(n14817), 
        .IN3(n10837), .IN4(\fadd_0_0_0_0_6/fracresultfar0 [6]), .IN5(
        \fadd_0_0_0_0_6/fracresultfar0 [4]), .IN6(
        \fadd_0_0_0_0_6/add_859/B[1] ), .Q(n10846) );
  AO222X1 U3644 ( .IN1(n10831), .IN2(n13699), .IN3(n10844), .IN4(n13563), 
        .IN5(n12844), .IN6(n10848), .Q(\fadd_0_0_0_0_6/resultbeforeround [2])
         );
  AO222X1 U3645 ( .IN1(\fadd_0_0_0_0_6/fracresultfar0 [4]), .IN2(n14817), 
        .IN3(\fadd_0_0_0_0_6/fracresultfar0 [5]), .IN4(n10837), .IN5(
        \fadd_0_0_0_0_6/add_859/B[1] ), .IN6(
        \fadd_0_0_0_0_6/fracresultfar0 [3]), .Q(n10848) );
  AO222X1 U3647 ( .IN1(n10831), .IN2(n13563), .IN3(n10844), .IN4(n13486), 
        .IN5(n12844), .IN6(n10849), .Q(\fadd_0_0_0_0_6/resultbeforeround [1])
         );
  AO222X1 U3648 ( .IN1(\fadd_0_0_0_0_6/fracresultfar0 [3]), .IN2(n14817), 
        .IN3(\fadd_0_0_0_0_6/fracresultfar0 [4]), .IN4(n10837), .IN5(
        \fadd_0_0_0_0_6/add_859/B[1] ), .IN6(
        \fadd_0_0_0_0_6/fracresultfar0 [2]), .Q(n10849) );
  AO22X1 U3650 ( .IN1(n13647), .IN2(\fadd_0_0_0_0_6/exponentresultclose_d1 [6]), .IN3(\fadd_0_0_0_0_6/exponentresultfar1 [6]), .IN4(n12844), .Q(
        \fadd_0_0_0_0_6/resultbeforeround [10]) );
  AO222X1 U3651 ( .IN1(n10831), .IN2(n13486), .IN3(n10844), .IN4(n13678), 
        .IN5(n12844), .IN6(n10839), .Q(\fadd_0_0_0_0_6/resultbeforeround [0])
         );
  AO222X1 U3652 ( .IN1(\fadd_0_0_0_0_6/fracresultfar0 [2]), .IN2(n14817), 
        .IN3(\fadd_0_0_0_0_6/fracresultfar0 [3]), .IN4(n10837), .IN5(
        \fadd_0_0_0_0_6/fracresultfar0 [1]), .IN6(
        \fadd_0_0_0_0_6/add_859/B[1] ), .Q(n10839) );
  AND2X1 U3659 ( .IN1(n12861), .IN2(n13647), .Q(n10831) );
  OA221X1 U3661 ( .IN1(n10850), .IN2(n10851), .IN3(n10852), .IN4(n10853), 
        .IN5(n10854), .Q(\fadd_0_0_0_0_6/ressign ) );
  XOR2X1 U3662 ( .IN1(n10855), .IN2(n10856), .Q(n10854) );
  OR3X1 U3663 ( .IN1(\fadd_0_0_0_0_6/fracrcloseymx [0]), .IN2(
        \fadd_0_0_0_0_6/fracrcloseymx [1]), .IN3(n10855), .Q(n10853) );
  OR4X1 U3666 ( .IN1(\fadd_0_0_0_0_6/fracrcloseymx [2]), .IN2(
        \fadd_0_0_0_0_6/fracrcloseymx [3]), .IN3(
        \fadd_0_0_0_0_6/fracrcloseymx [4]), .IN4(
        \fadd_0_0_0_0_6/fracrcloseymx [5]), .Q(n10852) );
  OR4X1 U3667 ( .IN1(n10857), .IN2(\fadd_0_0_0_0_6/fracrcloseymx [0]), .IN3(
        \fadd_0_0_0_0_6/fracrclosexmy [1]), .IN4(
        \fadd_0_0_0_0_6/fracrclosexmy [2]), .Q(n10851) );
  AO21X1 U3668 ( .IN1(n10858), .IN2(n10859), .IN3(n14805), .Q(n10857) );
  NAND4X0 U3669 ( .IN1(n10861), .IN2(n10862), .IN3(n14813), .IN4(n14812), .QN(
        n10859) );
  NAND4X0 U3670 ( .IN1(n10865), .IN2(n14309), .IN3(n14815), .IN4(n14814), .QN(
        n10858) );
  AO21X1 U3672 ( .IN1(\fadd_0_0_0_0_6/sub_784/B[1] ), .IN2(n14054), .IN3(
        n10870), .Q(\fadd_0_0_0_0_6/norm/level1 [4]) );
  OAI22X1 U3674 ( .IN1(n14934), .IN2(n11559), .IN3(n10871), .IN4(n11909), .QN(
        \fadd_0_0_0_0_6/norm/level1 [3]) );
  OAI22X1 U3675 ( .IN1(n14934), .IN2(n11558), .IN3(n10871), .IN4(n11910), .QN(
        \fadd_0_0_0_0_6/norm/level1 [2]) );
  NOR3X0 U3680 ( .IN1(n13542), .IN2(n8656), .IN3(n10870), .QN(
        \fadd_0_0_0_0_6/sub_784/B[1] ) );
  OAI21X1 U3681 ( .IN1(n10416), .IN2(n11558), .IN3(n11908), .QN(n10870) );
  NAND4X0 U3684 ( .IN1(n11907), .IN2(n11908), .IN3(n11909), .IN4(n11910), .QN(
        n10416) );
  AO22X1 U3685 ( .IN1(n14309), .IN2(n13508), .IN3(n10862), .IN4(n13471), .Q(
        \fadd_0_0_0_0_6/newy_11 ) );
  AO22X1 U3686 ( .IN1(n14309), .IN2(n13473), .IN3(n10862), .IN4(n13590), .Q(
        \fadd_0_0_0_0_6/newy_10 ) );
  AO22X1 U3687 ( .IN1(n14309), .IN2(n5554), .IN3(n10862), .IN4(n5566), .Q(
        \fadd_0_0_0_0_6/newx [8]) );
  AO22X1 U3690 ( .IN1(n14309), .IN2(n5553), .IN3(n10862), .IN4(n5565), .Q(
        \fadd_0_0_0_0_6/newx [7]) );
  AO22X1 U3693 ( .IN1(n14309), .IN2(n5552), .IN3(n10862), .IN4(n5564), .Q(
        \fadd_0_0_0_0_6/newx [6]) );
  AO22X1 U3696 ( .IN1(n14309), .IN2(n5551), .IN3(n10862), .IN4(n5563), .Q(
        \fadd_0_0_0_0_6/newx [5]) );
  AO22X1 U3699 ( .IN1(n14309), .IN2(n5550), .IN3(n10862), .IN4(n5562), .Q(
        \fadd_0_0_0_0_6/newx [4]) );
  AO22X1 U3702 ( .IN1(n14309), .IN2(n13578), .IN3(n10862), .IN4(n13496), .Q(
        \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ) );
  AO22X1 U3705 ( .IN1(n14309), .IN2(n13561), .IN3(n10862), .IN4(n13494), .Q(
        \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ) );
  AO22X1 U3708 ( .IN1(n14309), .IN2(n13536), .IN3(n10862), .IN4(n13481), .Q(
        \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ) );
  AO22X1 U3712 ( .IN1(n14309), .IN2(n13590), .IN3(n10862), .IN4(n13473), .Q(
        \fadd_0_0_0_0_6/newx [10]) );
  AO22X1 U3714 ( .IN1(n14309), .IN2(n13525), .IN3(n10862), .IN4(n13479), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ) );
  XOR2X1 U3717 ( .IN1(n10872), .IN2(n14805), .Q(
        \fadd_0_0_0_0_6/fracyfarxorop [6]) );
  XOR2X1 U3719 ( .IN1(n10875), .IN2(n12754), .Q(
        \fadd_0_0_0_0_6/fracyfarxorop [5]) );
  OA21X1 U3720 ( .IN1(n12751), .IN2(n14807), .IN3(n14802), .Q(n10875) );
  XOR2X1 U3722 ( .IN1(n10878), .IN2(n12754), .Q(
        \fadd_0_0_0_0_6/fracyfarxorop [4]) );
  OA22X1 U3723 ( .IN1(n14804), .IN2(n10879), .IN3(n12751), .IN4(n10880), .Q(
        n10878) );
  AO22X1 U3725 ( .IN1(n10882), .IN2(n14804), .IN3(n10883), .IN4(n12751), .Q(
        \fadd_0_0_0_0_6/fracyfarxorop [3]) );
  XOR2X1 U3726 ( .IN1(n10880), .IN2(n12754), .Q(n10883) );
  AO21X1 U3727 ( .IN1(n14808), .IN2(n10885), .IN3(n14801), .Q(n10880) );
  AO22X1 U3728 ( .IN1(n10887), .IN2(n14804), .IN3(n10882), .IN4(n12751), .Q(
        \fadd_0_0_0_0_6/fracyfarxorop [2]) );
  XOR2X1 U3729 ( .IN1(n14805), .IN2(n10888), .Q(n10882) );
  OA22X1 U3730 ( .IN1(n10881), .IN2(n10889), .IN3(n10890), .IN4(n10877), .Q(
        n10888) );
  AO22X1 U3732 ( .IN1(n10892), .IN2(n14804), .IN3(n10887), .IN4(n12751), .Q(
        \fadd_0_0_0_0_6/fracyfarxorop [1]) );
  XOR2X1 U3733 ( .IN1(n14805), .IN2(n10893), .Q(n10887) );
  OA22X1 U3734 ( .IN1(n10894), .IN2(n10889), .IN3(n14803), .IN4(n10895), .Q(
        n10893) );
  AO22X1 U3736 ( .IN1(n10892), .IN2(n12751), .IN3(n10896), .IN4(n14804), .Q(
        \fadd_0_0_0_0_6/fracyfarxorop [0]) );
  XOR2X1 U3738 ( .IN1(n12752), .IN2(n12754), .Q(n10896) );
  OA22X1 U3739 ( .IN1(n14803), .IN2(n12753), .IN3(n14810), .IN4(n14800), .Q(
        n12752) );
  XOR2X1 U3743 ( .IN1(n14805), .IN2(n10898), .Q(n10892) );
  AOI22X1 U3744 ( .IN1(n14809), .IN2(n14801), .IN3(n10891), .IN4(
        \fadd_0_0_0_0_6/rightshiftercomponent/level2[1] ), .QN(n10898) );
  OA221X1 U3748 ( .IN1(n14812), .IN2(n14309), .IN3(n14814), .IN4(n10862), 
        .IN5(n10897), .Q(n10885) );
  OA221X1 U3752 ( .IN1(n14813), .IN2(n14309), .IN3(n14815), .IN4(n10862), 
        .IN5(n10897), .Q(n10891) );
  OA22X1 U3753 ( .IN1(n14309), .IN2(n10861), .IN3(n10865), .IN4(n10862), .Q(
        n10897) );
  XOR2X1 U3759 ( .IN1(n14806), .IN2(\fadd_0_0_0_0_6/newy_9 ), .Q(n12754) );
  OAI22X1 U3760 ( .IN1(n10862), .IN2(n11781), .IN3(n14309), .IN4(n11770), .QN(
        \fadd_0_0_0_0_6/newy_9 ) );
  OA22X1 U3762 ( .IN1(n10862), .IN2(n11770), .IN3(n14309), .IN4(n11781), .Q(
        n10856) );
  AO22X1 U3764 ( .IN1(n14811), .IN2(n14808), .IN3(n14807), .IN4(n10899), .Q(
        \fadd_0_0_0_0_6/fracyclose1 [3]) );
  OA22X1 U3766 ( .IN1(n10862), .IN2(n11775), .IN3(n14309), .IN4(n11764), .Q(
        n10881) );
  AO22X1 U3767 ( .IN1(n14811), .IN2(n14809), .IN3(n14808), .IN4(n10899), .Q(
        \fadd_0_0_0_0_6/fracyclose1 [2]) );
  OA22X1 U3769 ( .IN1(n10862), .IN2(n11774), .IN3(n14309), .IN4(n11763), .Q(
        n10894) );
  AO22X1 U3770 ( .IN1(n14809), .IN2(n10899), .IN3(n14811), .IN4(n14810), .Q(
        \fadd_0_0_0_0_6/fracyclose1 [1]) );
  OA22X1 U3773 ( .IN1(n10862), .IN2(n11773), .IN3(n14309), .IN4(n11762), .Q(
        n10890) );
  OA22X1 U3775 ( .IN1(n10862), .IN2(n11772), .IN3(n14309), .IN4(n11761), .Q(
        n10900) );
  AO22X1 U3777 ( .IN1(\fadd_0_0_0_0_6/exponentdifferenceyx [0]), .IN2(n14309), 
        .IN3(\fadd_0_0_0_0_6/exponentdifferencexy [0]), .IN4(n10862), .Q(
        n10899) );
  OA22X1 U3780 ( .IN1(n11771), .IN2(n10903), .IN3(
        \fadd_0_0_0_0_6/sub_707/carry [5]), .IN4(n13473), .Q(n10902) );
  AO22X1 U3787 ( .IN1(\fadd_0_0_0_0_6/fracrcloseymx [5]), .IN2(n14115), .IN3(
        \fadd_0_0_0_0_6/fracrclosexmy [5]), .IN4(n14646), .Q(
        \fadd_0_0_0_0_6/fracrclose1 [5]) );
  AO22X1 U3788 ( .IN1(\fadd_0_0_0_0_6/fracrcloseymx [4]), .IN2(n14115), .IN3(
        \fadd_0_0_0_0_6/fracrclosexmy [4]), .IN4(n14646), .Q(
        \fadd_0_0_0_0_6/fracrclose1 [4]) );
  AO22X1 U3789 ( .IN1(\fadd_0_0_0_0_6/fracrcloseymx [3]), .IN2(n14115), .IN3(
        \fadd_0_0_0_0_6/fracrclosexmy [3]), .IN4(n14646), .Q(
        \fadd_0_0_0_0_6/fracrclose1 [3]) );
  AO22X1 U3790 ( .IN1(\fadd_0_0_0_0_6/fracrcloseymx [2]), .IN2(n14115), .IN3(
        \fadd_0_0_0_0_6/fracrclosexmy [2]), .IN4(n14646), .Q(
        \fadd_0_0_0_0_6/fracrclose1 [2]) );
  AO22X1 U3791 ( .IN1(\fadd_0_0_0_0_6/fracrcloseymx [1]), .IN2(n14115), .IN3(
        \fadd_0_0_0_0_6/fracrclosexmy [1]), .IN4(n14646), .Q(
        \fadd_0_0_0_0_6/fracrclose1 [1]) );
  AO22X1 U3792 ( .IN1(\fadd_0_0_0_0_6/fracrcloseymx [0]), .IN2(n14115), .IN3(
        \fadd_0_0_0_0_6/fracrcloseymx [0]), .IN4(n14646), .Q(
        \fadd_0_0_0_0_6/fracrclose1 [0]) );
  NOR3X0 U3796 ( .IN1(n14953), .IN2(n11557), .IN3(n10838), .QN(
        \fadd_0_0_0_0_6/cinaddfar ) );
  AND2X1 U3797 ( .IN1(\fadd_0_0_0_0_6/rightshiftercomponent/level1_d2[0] ), 
        .IN2(\fadd_0_0_0_0_6/rightshiftercomponent/ps_d2[0] ), .Q(n10838) );
  NOR3X0 U3799 ( .IN1(n14933), .IN2(n11555), .IN3(n10415), .QN(
        \fadd_0_0_0_0_5/zerofromclose ) );
  NAND3X0 U3801 ( .IN1(n13682), .IN2(n13490), .IN3(n10912), .QN(n10909) );
  NAND3X0 U3802 ( .IN1(n10913), .IN2(n10914), .IN3(n12843), .QN(n10908) );
  AO222X1 U3807 ( .IN1(\fadd_0_0_0_0_5/fracresultfar0 [1]), .IN2(n14796), 
        .IN3(\fadd_0_0_0_0_5/fracresultfar0 [2]), .IN4(n10918), .IN5(
        \fadd_0_0_0_0_5/fracresultfar0 [0]), .IN6(n14229), .Q(n10913) );
  AO22X1 U3808 ( .IN1(n10922), .IN2(
        \fadd_0_0_0_0_5/rightshiftercomponent/ps_d1 [1]), .IN3(n10923), .IN4(
        \fadd_0_0_0_0_5/rightshiftercomponent/ps_d1 [2]), .Q(
        \fadd_0_0_0_0_5/rightshiftercomponent/n389_o ) );
  AO22X1 U3811 ( .IN1(n13651), .IN2(\fadd_0_0_0_0_5/exponentresultclose_d1 [5]), .IN3(\fadd_0_0_0_0_5/exponentresultfar1 [5]), .IN4(n12843), .Q(
        \fadd_0_0_0_0_5/resultbeforeround [9]) );
  AO22X1 U3812 ( .IN1(n13651), .IN2(\fadd_0_0_0_0_5/exponentresultclose_d1 [4]), .IN3(\fadd_0_0_0_0_5/exponentresultfar1 [4]), .IN4(n12843), .Q(
        \fadd_0_0_0_0_5/resultbeforeround [8]) );
  AO22X1 U3813 ( .IN1(n13651), .IN2(\fadd_0_0_0_0_5/exponentresultclose_d1 [3]), .IN3(\fadd_0_0_0_0_5/exponentresultfar1 [3]), .IN4(n12843), .Q(
        \fadd_0_0_0_0_5/resultbeforeround [7]) );
  AO22X1 U3814 ( .IN1(n13651), .IN2(\fadd_0_0_0_0_5/exponentresultclose_d1 [2]), .IN3(\fadd_0_0_0_0_5/exponentresultfar1 [2]), .IN4(n12843), .Q(
        \fadd_0_0_0_0_5/resultbeforeround [6]) );
  AO22X1 U3815 ( .IN1(n13651), .IN2(\fadd_0_0_0_0_5/exponentresultclose_d1 [1]), .IN3(\fadd_0_0_0_0_5/exponentresultfar1 [1]), .IN4(n12843), .Q(
        \fadd_0_0_0_0_5/resultbeforeround [5]) );
  AO22X1 U3816 ( .IN1(n13651), .IN2(\fadd_0_0_0_0_5/exponentresultclose_d1 [0]), .IN3(\fadd_0_0_0_0_5/exponentresultfar1 [0]), .IN4(n12843), .Q(
        \fadd_0_0_0_0_5/resultbeforeround [4]) );
  AO222X1 U3817 ( .IN1(n10912), .IN2(\fadd_0_0_0_0_5/norm/level1_d1[4] ), 
        .IN3(n10925), .IN4(n13703), .IN5(n12843), .IN6(n10927), .Q(
        \fadd_0_0_0_0_5/resultbeforeround [3]) );
  AO222X1 U3818 ( .IN1(\fadd_0_0_0_0_5/fracresultfar0 [5]), .IN2(n14796), 
        .IN3(n10918), .IN4(\fadd_0_0_0_0_5/fracresultfar0 [6]), .IN5(
        \fadd_0_0_0_0_5/fracresultfar0 [4]), .IN6(n14229), .Q(n10927) );
  AO222X1 U3819 ( .IN1(n10912), .IN2(n13703), .IN3(n10925), .IN4(n13567), 
        .IN5(n12843), .IN6(n10929), .Q(\fadd_0_0_0_0_5/resultbeforeround [2])
         );
  AO222X1 U3820 ( .IN1(\fadd_0_0_0_0_5/fracresultfar0 [4]), .IN2(n14796), 
        .IN3(\fadd_0_0_0_0_5/fracresultfar0 [5]), .IN4(n10918), .IN5(n14229), 
        .IN6(\fadd_0_0_0_0_5/fracresultfar0 [3]), .Q(n10929) );
  AO222X1 U3822 ( .IN1(n10912), .IN2(n13567), .IN3(n10925), .IN4(n13490), 
        .IN5(n12843), .IN6(n10930), .Q(\fadd_0_0_0_0_5/resultbeforeround [1])
         );
  AO222X1 U3823 ( .IN1(\fadd_0_0_0_0_5/fracresultfar0 [3]), .IN2(n14796), 
        .IN3(\fadd_0_0_0_0_5/fracresultfar0 [4]), .IN4(n10918), .IN5(n14229), 
        .IN6(\fadd_0_0_0_0_5/fracresultfar0 [2]), .Q(n10930) );
  AO22X1 U3825 ( .IN1(n13651), .IN2(\fadd_0_0_0_0_5/exponentresultclose_d1 [6]), .IN3(\fadd_0_0_0_0_5/exponentresultfar1 [6]), .IN4(n12843), .Q(
        \fadd_0_0_0_0_5/resultbeforeround [10]) );
  AO222X1 U3826 ( .IN1(n10912), .IN2(n13490), .IN3(n10925), .IN4(n13682), 
        .IN5(n12843), .IN6(n10920), .Q(\fadd_0_0_0_0_5/resultbeforeround [0])
         );
  AO222X1 U3827 ( .IN1(\fadd_0_0_0_0_5/fracresultfar0 [2]), .IN2(n14796), 
        .IN3(\fadd_0_0_0_0_5/fracresultfar0 [3]), .IN4(n10918), .IN5(
        \fadd_0_0_0_0_5/fracresultfar0 [1]), .IN6(n14229), .Q(n10920) );
  AND2X1 U3834 ( .IN1(n12859), .IN2(n13651), .Q(n10912) );
  OA221X1 U3836 ( .IN1(n10931), .IN2(n10932), .IN3(n10933), .IN4(n10934), 
        .IN5(n10935), .Q(\fadd_0_0_0_0_5/ressign ) );
  OR4X1 U3841 ( .IN1(\fadd_0_0_0_0_5/fracrcloseymx [2]), .IN2(
        \fadd_0_0_0_0_5/fracrcloseymx [3]), .IN3(
        \fadd_0_0_0_0_5/fracrcloseymx [4]), .IN4(
        \fadd_0_0_0_0_5/fracrcloseymx [5]), .Q(n10933) );
  OR4X1 U3842 ( .IN1(n10938), .IN2(\fadd_0_0_0_0_5/fracrcloseymx [0]), .IN3(
        \fadd_0_0_0_0_5/fracrclosexmy [1]), .IN4(
        \fadd_0_0_0_0_5/fracrclosexmy [2]), .Q(n10932) );
  AO21X1 U3843 ( .IN1(n10939), .IN2(n10940), .IN3(n14784), .Q(n10938) );
  NAND4X0 U3844 ( .IN1(n10942), .IN2(n10943), .IN3(n14792), .IN4(n14791), .QN(
        n10940) );
  NAND4X0 U3845 ( .IN1(n10946), .IN2(n14308), .IN3(n14794), .IN4(n14793), .QN(
        n10939) );
  AO21X1 U3847 ( .IN1(\fadd_0_0_0_0_5/sub_784/B[1] ), .IN2(n14053), .IN3(
        n10951), .Q(\fadd_0_0_0_0_5/norm/level1 [4]) );
  OAI22X1 U3849 ( .IN1(n14933), .IN2(n11546), .IN3(n10952), .IN4(n11905), .QN(
        \fadd_0_0_0_0_5/norm/level1 [3]) );
  OAI22X1 U3850 ( .IN1(n14933), .IN2(n11545), .IN3(n10952), .IN4(n11906), .QN(
        \fadd_0_0_0_0_5/norm/level1 [2]) );
  NOR3X0 U3855 ( .IN1(n13543), .IN2(n8652), .IN3(n10951), .QN(
        \fadd_0_0_0_0_5/sub_784/B[1] ) );
  OAI21X1 U3856 ( .IN1(n10415), .IN2(n11545), .IN3(n11904), .QN(n10951) );
  NAND4X0 U3859 ( .IN1(n11903), .IN2(n11904), .IN3(n11905), .IN4(n11906), .QN(
        n10415) );
  AO22X1 U3860 ( .IN1(n14308), .IN2(n13511), .IN3(n10943), .IN4(n13624), .Q(
        \fadd_0_0_0_0_5/newy_11 ) );
  AO22X1 U3861 ( .IN1(n14308), .IN2(n13503), .IN3(n10943), .IN4(n13891), .Q(
        \fadd_0_0_0_0_5/newy_10 ) );
  AO22X1 U3862 ( .IN1(n14308), .IN2(n5626), .IN3(n10943), .IN4(n5638), .Q(
        \fadd_0_0_0_0_5/newx [8]) );
  AO22X1 U3865 ( .IN1(n14308), .IN2(n5625), .IN3(n10943), .IN4(n5637), .Q(
        \fadd_0_0_0_0_5/newx [7]) );
  AO22X1 U3868 ( .IN1(n14308), .IN2(n5624), .IN3(n10943), .IN4(n5636), .Q(
        \fadd_0_0_0_0_5/newx [6]) );
  AO22X1 U3871 ( .IN1(n14308), .IN2(n5623), .IN3(n10943), .IN4(n5635), .Q(
        \fadd_0_0_0_0_5/newx [5]) );
  AO22X1 U3874 ( .IN1(n14308), .IN2(n5622), .IN3(n10943), .IN4(n5634), .Q(
        \fadd_0_0_0_0_5/newx [4]) );
  AO22X1 U3877 ( .IN1(n14308), .IN2(n13710), .IN3(n10943), .IN4(n13572), .Q(
        \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ) );
  AO22X1 U3880 ( .IN1(n14308), .IN2(n13688), .IN3(n10943), .IN4(n13555), .Q(
        \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ) );
  AO22X1 U3883 ( .IN1(n14308), .IN2(n13667), .IN3(n10943), .IN4(n13530), .Q(
        \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ) );
  AO22X1 U3887 ( .IN1(n14308), .IN2(n13891), .IN3(n10943), .IN4(n13503), .Q(
        \fadd_0_0_0_0_5/newx [10]) );
  AO22X1 U3889 ( .IN1(n14308), .IN2(n13639), .IN3(n10943), .IN4(n13519), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ) );
  XOR2X1 U3892 ( .IN1(n10953), .IN2(n14784), .Q(
        \fadd_0_0_0_0_5/fracyfarxorop [6]) );
  XOR2X1 U3894 ( .IN1(n10956), .IN2(n12742), .Q(
        \fadd_0_0_0_0_5/fracyfarxorop [5]) );
  OA21X1 U3895 ( .IN1(n12739), .IN2(n14786), .IN3(n14781), .Q(n10956) );
  XOR2X1 U3897 ( .IN1(n10959), .IN2(n12742), .Q(
        \fadd_0_0_0_0_5/fracyfarxorop [4]) );
  OA22X1 U3898 ( .IN1(n14783), .IN2(n10960), .IN3(n12739), .IN4(n10961), .Q(
        n10959) );
  AO22X1 U3900 ( .IN1(n10963), .IN2(n14783), .IN3(n10964), .IN4(n12739), .Q(
        \fadd_0_0_0_0_5/fracyfarxorop [3]) );
  XOR2X1 U3901 ( .IN1(n10961), .IN2(n12742), .Q(n10964) );
  AO21X1 U3902 ( .IN1(n14787), .IN2(n10966), .IN3(n14780), .Q(n10961) );
  AO22X1 U3903 ( .IN1(n10968), .IN2(n14783), .IN3(n10963), .IN4(n12739), .Q(
        \fadd_0_0_0_0_5/fracyfarxorop [2]) );
  XOR2X1 U3904 ( .IN1(n14784), .IN2(n10969), .Q(n10963) );
  OA22X1 U3905 ( .IN1(n10962), .IN2(n10970), .IN3(n10971), .IN4(n10958), .Q(
        n10969) );
  AO22X1 U3907 ( .IN1(n10973), .IN2(n14783), .IN3(n10968), .IN4(n12739), .Q(
        \fadd_0_0_0_0_5/fracyfarxorop [1]) );
  XOR2X1 U3908 ( .IN1(n14784), .IN2(n10974), .Q(n10968) );
  OA22X1 U3909 ( .IN1(n10975), .IN2(n10970), .IN3(n14782), .IN4(n10976), .Q(
        n10974) );
  AO22X1 U3911 ( .IN1(n10973), .IN2(n12739), .IN3(n10977), .IN4(n14783), .Q(
        \fadd_0_0_0_0_5/fracyfarxorop [0]) );
  XOR2X1 U3913 ( .IN1(n12740), .IN2(n12742), .Q(n10977) );
  OA22X1 U3914 ( .IN1(n14782), .IN2(n12741), .IN3(n14789), .IN4(n14779), .Q(
        n12740) );
  XOR2X1 U3918 ( .IN1(n14784), .IN2(n10979), .Q(n10973) );
  AOI22X1 U3919 ( .IN1(n14788), .IN2(n14780), .IN3(n10972), .IN4(
        \fadd_0_0_0_0_5/rightshiftercomponent/level2[1] ), .QN(n10979) );
  OA221X1 U3923 ( .IN1(n14791), .IN2(n14308), .IN3(n14793), .IN4(n10943), 
        .IN5(n10978), .Q(n10966) );
  OA221X1 U3927 ( .IN1(n14792), .IN2(n14308), .IN3(n14794), .IN4(n10943), 
        .IN5(n10978), .Q(n10972) );
  OA22X1 U3928 ( .IN1(n14308), .IN2(n10942), .IN3(n10946), .IN4(n10943), .Q(
        n10978) );
  XOR2X1 U3934 ( .IN1(n14785), .IN2(\fadd_0_0_0_0_5/newy_9 ), .Q(n12742) );
  AO22X1 U3935 ( .IN1(n14308), .IN2(n13581), .IN3(n10943), .IN4(n13719), .Q(
        \fadd_0_0_0_0_5/newy_9 ) );
  OA22X1 U3939 ( .IN1(n10943), .IN2(n11728), .IN3(n14308), .IN4(n11739), .Q(
        n10937) );
  AO22X1 U3941 ( .IN1(n14790), .IN2(n14787), .IN3(n14786), .IN4(n10980), .Q(
        \fadd_0_0_0_0_5/fracyclose1 [3]) );
  OA22X1 U3943 ( .IN1(n10943), .IN2(n11733), .IN3(n14308), .IN4(n11722), .Q(
        n10962) );
  AO22X1 U3944 ( .IN1(n14790), .IN2(n14788), .IN3(n14787), .IN4(n10980), .Q(
        \fadd_0_0_0_0_5/fracyclose1 [2]) );
  OA22X1 U3946 ( .IN1(n10943), .IN2(n11732), .IN3(n14308), .IN4(n11721), .Q(
        n10975) );
  AO22X1 U3947 ( .IN1(n14788), .IN2(n10980), .IN3(n14790), .IN4(n14789), .Q(
        \fadd_0_0_0_0_5/fracyclose1 [1]) );
  OA22X1 U3950 ( .IN1(n10943), .IN2(n11731), .IN3(n14308), .IN4(n11720), .Q(
        n10971) );
  OA22X1 U3952 ( .IN1(n10943), .IN2(n11730), .IN3(n14308), .IN4(n11719), .Q(
        n10981) );
  AO22X1 U3954 ( .IN1(\fadd_0_0_0_0_5/exponentdifferenceyx [0]), .IN2(n14308), 
        .IN3(\fadd_0_0_0_0_5/exponentdifferencexy [0]), .IN4(n10943), .Q(
        n10980) );
  OA22X1 U3957 ( .IN1(n11729), .IN2(n10984), .IN3(
        \fadd_0_0_0_0_5/sub_707/carry [5]), .IN4(n13503), .Q(n10983) );
  AO22X1 U3964 ( .IN1(\fadd_0_0_0_0_5/fracrcloseymx [5]), .IN2(n14111), .IN3(
        \fadd_0_0_0_0_5/fracrclosexmy [5]), .IN4(n14644), .Q(
        \fadd_0_0_0_0_5/fracrclose1 [5]) );
  AO22X1 U3965 ( .IN1(\fadd_0_0_0_0_5/fracrcloseymx [4]), .IN2(n14111), .IN3(
        \fadd_0_0_0_0_5/fracrclosexmy [4]), .IN4(n14644), .Q(
        \fadd_0_0_0_0_5/fracrclose1 [4]) );
  AO22X1 U3966 ( .IN1(\fadd_0_0_0_0_5/fracrcloseymx [3]), .IN2(n14111), .IN3(
        \fadd_0_0_0_0_5/fracrclosexmy [3]), .IN4(n14644), .Q(
        \fadd_0_0_0_0_5/fracrclose1 [3]) );
  AO22X1 U3967 ( .IN1(\fadd_0_0_0_0_5/fracrcloseymx [2]), .IN2(n14111), .IN3(
        \fadd_0_0_0_0_5/fracrclosexmy [2]), .IN4(n14644), .Q(
        \fadd_0_0_0_0_5/fracrclose1 [2]) );
  AO22X1 U3968 ( .IN1(\fadd_0_0_0_0_5/fracrcloseymx [1]), .IN2(n14111), .IN3(
        \fadd_0_0_0_0_5/fracrclosexmy [1]), .IN4(n14644), .Q(
        \fadd_0_0_0_0_5/fracrclose1 [1]) );
  AO22X1 U3969 ( .IN1(\fadd_0_0_0_0_5/fracrcloseymx [0]), .IN2(n14111), .IN3(
        \fadd_0_0_0_0_5/fracrcloseymx [0]), .IN4(n14644), .Q(
        \fadd_0_0_0_0_5/fracrclose1 [0]) );
  NOR3X0 U3973 ( .IN1(n14949), .IN2(n11544), .IN3(n10919), .QN(
        \fadd_0_0_0_0_5/cinaddfar ) );
  AND2X1 U3974 ( .IN1(\fadd_0_0_0_0_5/rightshiftercomponent/level1_d2[0] ), 
        .IN2(\fadd_0_0_0_0_5/rightshiftercomponent/ps_d2[0] ), .Q(n10919) );
  NOR3X0 U3976 ( .IN1(n14932), .IN2(n11542), .IN3(n10414), .QN(
        \fadd_0_0_0_0_4/zerofromclose ) );
  NAND3X0 U3978 ( .IN1(n13672), .IN2(n13483), .IN3(n10993), .QN(n10990) );
  NAND3X0 U3979 ( .IN1(n10994), .IN2(n10995), .IN3(n12842), .QN(n10989) );
  AO222X1 U3984 ( .IN1(\fadd_0_0_0_0_4/fracresultfar0 [1]), .IN2(n14775), 
        .IN3(\fadd_0_0_0_0_4/fracresultfar0 [2]), .IN4(n10999), .IN5(
        \fadd_0_0_0_0_4/fracresultfar0 [0]), .IN6(n14228), .Q(n10994) );
  AO22X1 U3985 ( .IN1(n11003), .IN2(
        \fadd_0_0_0_0_4/rightshiftercomponent/ps_d1 [1]), .IN3(n11004), .IN4(
        \fadd_0_0_0_0_4/rightshiftercomponent/ps_d1 [2]), .Q(
        \fadd_0_0_0_0_4/rightshiftercomponent/n389_o ) );
  AO22X1 U3988 ( .IN1(n13644), .IN2(\fadd_0_0_0_0_4/exponentresultclose_d1 [5]), .IN3(\fadd_0_0_0_0_4/exponentresultfar1 [5]), .IN4(n12842), .Q(
        \fadd_0_0_0_0_4/resultbeforeround [9]) );
  AO22X1 U3989 ( .IN1(n13644), .IN2(\fadd_0_0_0_0_4/exponentresultclose_d1 [4]), .IN3(\fadd_0_0_0_0_4/exponentresultfar1 [4]), .IN4(n12842), .Q(
        \fadd_0_0_0_0_4/resultbeforeround [8]) );
  AO22X1 U3990 ( .IN1(n13644), .IN2(\fadd_0_0_0_0_4/exponentresultclose_d1 [3]), .IN3(\fadd_0_0_0_0_4/exponentresultfar1 [3]), .IN4(n12842), .Q(
        \fadd_0_0_0_0_4/resultbeforeround [7]) );
  AO22X1 U3991 ( .IN1(n13644), .IN2(\fadd_0_0_0_0_4/exponentresultclose_d1 [2]), .IN3(\fadd_0_0_0_0_4/exponentresultfar1 [2]), .IN4(n12842), .Q(
        \fadd_0_0_0_0_4/resultbeforeround [6]) );
  AO22X1 U3992 ( .IN1(n13644), .IN2(\fadd_0_0_0_0_4/exponentresultclose_d1 [1]), .IN3(\fadd_0_0_0_0_4/exponentresultfar1 [1]), .IN4(n12842), .Q(
        \fadd_0_0_0_0_4/resultbeforeround [5]) );
  AO22X1 U3993 ( .IN1(n13644), .IN2(\fadd_0_0_0_0_4/exponentresultclose_d1 [0]), .IN3(\fadd_0_0_0_0_4/exponentresultfar1 [0]), .IN4(n12842), .Q(
        \fadd_0_0_0_0_4/resultbeforeround [4]) );
  AO222X1 U3994 ( .IN1(n10993), .IN2(\fadd_0_0_0_0_4/norm/level1_d1[4] ), 
        .IN3(n11006), .IN4(n13693), .IN5(n12842), .IN6(n11008), .Q(
        \fadd_0_0_0_0_4/resultbeforeround [3]) );
  AO222X1 U3995 ( .IN1(\fadd_0_0_0_0_4/fracresultfar0 [5]), .IN2(n14775), 
        .IN3(n10999), .IN4(\fadd_0_0_0_0_4/fracresultfar0 [6]), .IN5(
        \fadd_0_0_0_0_4/fracresultfar0 [4]), .IN6(n14228), .Q(n11008) );
  AO222X1 U3996 ( .IN1(n10993), .IN2(n13693), .IN3(n11006), .IN4(n13551), 
        .IN5(n12842), .IN6(n11010), .Q(\fadd_0_0_0_0_4/resultbeforeround [2])
         );
  AO222X1 U3997 ( .IN1(\fadd_0_0_0_0_4/fracresultfar0 [4]), .IN2(n14775), 
        .IN3(\fadd_0_0_0_0_4/fracresultfar0 [5]), .IN4(n10999), .IN5(n14228), 
        .IN6(\fadd_0_0_0_0_4/fracresultfar0 [3]), .Q(n11010) );
  AO222X1 U3999 ( .IN1(n10993), .IN2(n13551), .IN3(n11006), .IN4(n13483), 
        .IN5(n12842), .IN6(n11011), .Q(\fadd_0_0_0_0_4/resultbeforeround [1])
         );
  AO222X1 U4000 ( .IN1(\fadd_0_0_0_0_4/fracresultfar0 [3]), .IN2(n14775), 
        .IN3(\fadd_0_0_0_0_4/fracresultfar0 [4]), .IN4(n10999), .IN5(n14228), 
        .IN6(\fadd_0_0_0_0_4/fracresultfar0 [2]), .Q(n11011) );
  AO22X1 U4002 ( .IN1(n13644), .IN2(\fadd_0_0_0_0_4/exponentresultclose_d1 [6]), .IN3(\fadd_0_0_0_0_4/exponentresultfar1 [6]), .IN4(n12842), .Q(
        \fadd_0_0_0_0_4/resultbeforeround [10]) );
  AO222X1 U4003 ( .IN1(n10993), .IN2(n13483), .IN3(n11006), .IN4(n13672), 
        .IN5(n12842), .IN6(n11001), .Q(\fadd_0_0_0_0_4/resultbeforeround [0])
         );
  AO222X1 U4004 ( .IN1(\fadd_0_0_0_0_4/fracresultfar0 [2]), .IN2(n14775), 
        .IN3(\fadd_0_0_0_0_4/fracresultfar0 [3]), .IN4(n10999), .IN5(
        \fadd_0_0_0_0_4/fracresultfar0 [1]), .IN6(n14228), .Q(n11001) );
  AND2X1 U4011 ( .IN1(n12857), .IN2(n13644), .Q(n10993) );
  OA221X1 U4013 ( .IN1(n11012), .IN2(n11013), .IN3(n11014), .IN4(n11015), 
        .IN5(n11016), .Q(\fadd_0_0_0_0_4/ressign ) );
  OR4X1 U4018 ( .IN1(\fadd_0_0_0_0_4/fracrcloseymx [2]), .IN2(
        \fadd_0_0_0_0_4/fracrcloseymx [3]), .IN3(
        \fadd_0_0_0_0_4/fracrcloseymx [4]), .IN4(
        \fadd_0_0_0_0_4/fracrcloseymx [5]), .Q(n11014) );
  OR4X1 U4019 ( .IN1(n11019), .IN2(\fadd_0_0_0_0_4/fracrcloseymx [0]), .IN3(
        \fadd_0_0_0_0_4/fracrclosexmy [1]), .IN4(
        \fadd_0_0_0_0_4/fracrclosexmy [2]), .Q(n11013) );
  AO21X1 U4020 ( .IN1(n11020), .IN2(n11021), .IN3(n14752), .Q(n11019) );
  NAND4X0 U4021 ( .IN1(n11023), .IN2(n11024), .IN3(n14760), .IN4(n14759), .QN(
        n11021) );
  NAND4X0 U4022 ( .IN1(n11027), .IN2(n14307), .IN3(n14762), .IN4(n14761), .QN(
        n11020) );
  AO21X1 U4024 ( .IN1(\fadd_0_0_0_0_4/sub_784/B[1] ), .IN2(n14052), .IN3(
        n11032), .Q(\fadd_0_0_0_0_4/norm/level1 [4]) );
  OAI22X1 U4026 ( .IN1(n14932), .IN2(n11533), .IN3(n11033), .IN4(n11901), .QN(
        \fadd_0_0_0_0_4/norm/level1 [3]) );
  OAI22X1 U4027 ( .IN1(n14932), .IN2(n11532), .IN3(n11033), .IN4(n11902), .QN(
        \fadd_0_0_0_0_4/norm/level1 [2]) );
  NOR3X0 U4032 ( .IN1(n13544), .IN2(n8648), .IN3(n11032), .QN(
        \fadd_0_0_0_0_4/sub_784/B[1] ) );
  OAI21X1 U4033 ( .IN1(n10414), .IN2(n11532), .IN3(n11900), .QN(n11032) );
  NAND4X0 U4036 ( .IN1(n11899), .IN2(n11900), .IN3(n11901), .IN4(n11902), .QN(
        n10414) );
  AO22X1 U4037 ( .IN1(n14307), .IN2(n13514), .IN3(n11024), .IN4(n13621), .Q(
        \fadd_0_0_0_0_4/newy_11 ) );
  AO22X1 U4038 ( .IN1(n14307), .IN2(n13505), .IN3(n11024), .IN4(n13888), .Q(
        \fadd_0_0_0_0_4/newy_10 ) );
  AO22X1 U4039 ( .IN1(n14307), .IN2(n5698), .IN3(n11024), .IN4(n5710), .Q(
        \fadd_0_0_0_0_4/newx [8]) );
  AO22X1 U4042 ( .IN1(n14307), .IN2(n5697), .IN3(n11024), .IN4(n5709), .Q(
        \fadd_0_0_0_0_4/newx [7]) );
  AO22X1 U4045 ( .IN1(n14307), .IN2(n5696), .IN3(n11024), .IN4(n5708), .Q(
        \fadd_0_0_0_0_4/newx [6]) );
  AO22X1 U4048 ( .IN1(n14307), .IN2(n5695), .IN3(n11024), .IN4(n5707), .Q(
        \fadd_0_0_0_0_4/newx [5]) );
  AO22X1 U4051 ( .IN1(n14307), .IN2(n5694), .IN3(n11024), .IN4(n5706), .Q(
        \fadd_0_0_0_0_4/newx [4]) );
  AO22X1 U4054 ( .IN1(n14307), .IN2(n13707), .IN3(n11024), .IN4(n13575), .Q(
        \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ) );
  AO22X1 U4057 ( .IN1(n14307), .IN2(n13685), .IN3(n11024), .IN4(n13558), .Q(
        \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ) );
  AO22X1 U4060 ( .IN1(n14307), .IN2(n13664), .IN3(n11024), .IN4(n13533), .Q(
        \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ) );
  AO22X1 U4064 ( .IN1(n14307), .IN2(n13888), .IN3(n11024), .IN4(n13505), .Q(
        \fadd_0_0_0_0_4/newx [10]) );
  AO22X1 U4066 ( .IN1(n14307), .IN2(n13636), .IN3(n11024), .IN4(n13522), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ) );
  XOR2X1 U4069 ( .IN1(n11034), .IN2(n14752), .Q(
        \fadd_0_0_0_0_4/fracyfarxorop [6]) );
  XOR2X1 U4071 ( .IN1(n11037), .IN2(n12734), .Q(
        \fadd_0_0_0_0_4/fracyfarxorop [5]) );
  OA21X1 U4072 ( .IN1(n12731), .IN2(n14754), .IN3(n14749), .Q(n11037) );
  XOR2X1 U4074 ( .IN1(n11040), .IN2(n12734), .Q(
        \fadd_0_0_0_0_4/fracyfarxorop [4]) );
  OA22X1 U4075 ( .IN1(n14751), .IN2(n11041), .IN3(n12731), .IN4(n11042), .Q(
        n11040) );
  AO22X1 U4077 ( .IN1(n11044), .IN2(n14751), .IN3(n11045), .IN4(n12731), .Q(
        \fadd_0_0_0_0_4/fracyfarxorop [3]) );
  XOR2X1 U4078 ( .IN1(n11042), .IN2(n12734), .Q(n11045) );
  AO21X1 U4079 ( .IN1(n14755), .IN2(n11047), .IN3(n14748), .Q(n11042) );
  AO22X1 U4080 ( .IN1(n11049), .IN2(n14751), .IN3(n11044), .IN4(n12731), .Q(
        \fadd_0_0_0_0_4/fracyfarxorop [2]) );
  XOR2X1 U4081 ( .IN1(n14752), .IN2(n11050), .Q(n11044) );
  OA22X1 U4082 ( .IN1(n11043), .IN2(n11051), .IN3(n11052), .IN4(n11039), .Q(
        n11050) );
  AO22X1 U4084 ( .IN1(n11054), .IN2(n14751), .IN3(n11049), .IN4(n12731), .Q(
        \fadd_0_0_0_0_4/fracyfarxorop [1]) );
  XOR2X1 U4085 ( .IN1(n14752), .IN2(n11055), .Q(n11049) );
  OA22X1 U4086 ( .IN1(n11056), .IN2(n11051), .IN3(n14750), .IN4(n11057), .Q(
        n11055) );
  AO22X1 U4088 ( .IN1(n11054), .IN2(n12731), .IN3(n11058), .IN4(n14751), .Q(
        \fadd_0_0_0_0_4/fracyfarxorop [0]) );
  XOR2X1 U4090 ( .IN1(n12732), .IN2(n12734), .Q(n11058) );
  OA22X1 U4091 ( .IN1(n14750), .IN2(n12733), .IN3(n14757), .IN4(n14747), .Q(
        n12732) );
  XOR2X1 U4095 ( .IN1(n14752), .IN2(n11060), .Q(n11054) );
  AOI22X1 U4096 ( .IN1(n14756), .IN2(n14748), .IN3(n11053), .IN4(
        \fadd_0_0_0_0_4/rightshiftercomponent/level2[1] ), .QN(n11060) );
  OA221X1 U4100 ( .IN1(n14759), .IN2(n14307), .IN3(n14761), .IN4(n11024), 
        .IN5(n11059), .Q(n11047) );
  OA221X1 U4104 ( .IN1(n14760), .IN2(n14307), .IN3(n14762), .IN4(n11024), 
        .IN5(n11059), .Q(n11053) );
  OA22X1 U4105 ( .IN1(n14307), .IN2(n11023), .IN3(n11027), .IN4(n11024), .Q(
        n11059) );
  XOR2X1 U4111 ( .IN1(n14753), .IN2(\fadd_0_0_0_0_4/newy_9 ), .Q(n12734) );
  AO22X1 U4112 ( .IN1(n14307), .IN2(n13584), .IN3(n11024), .IN4(n13716), .Q(
        \fadd_0_0_0_0_4/newy_9 ) );
  OA22X1 U4116 ( .IN1(n11024), .IN2(n11791), .IN3(n14307), .IN4(n11802), .Q(
        n11018) );
  AO22X1 U4118 ( .IN1(n14758), .IN2(n14755), .IN3(n14754), .IN4(n11061), .Q(
        \fadd_0_0_0_0_4/fracyclose1 [3]) );
  OA22X1 U4120 ( .IN1(n11024), .IN2(n11796), .IN3(n14307), .IN4(n11785), .Q(
        n11043) );
  AO22X1 U4121 ( .IN1(n14758), .IN2(n14756), .IN3(n14755), .IN4(n11061), .Q(
        \fadd_0_0_0_0_4/fracyclose1 [2]) );
  OA22X1 U4123 ( .IN1(n11024), .IN2(n11795), .IN3(n14307), .IN4(n11784), .Q(
        n11056) );
  AO22X1 U4124 ( .IN1(n14756), .IN2(n11061), .IN3(n14758), .IN4(n14757), .Q(
        \fadd_0_0_0_0_4/fracyclose1 [1]) );
  OA22X1 U4127 ( .IN1(n11024), .IN2(n11794), .IN3(n14307), .IN4(n11783), .Q(
        n11052) );
  OA22X1 U4129 ( .IN1(n11024), .IN2(n11793), .IN3(n14307), .IN4(n11782), .Q(
        n11062) );
  AO22X1 U4131 ( .IN1(\fadd_0_0_0_0_4/exponentdifferenceyx [0]), .IN2(n14307), 
        .IN3(\fadd_0_0_0_0_4/exponentdifferencexy [0]), .IN4(n11024), .Q(
        n11061) );
  OA22X1 U4134 ( .IN1(n11792), .IN2(n11065), .IN3(
        \fadd_0_0_0_0_4/sub_707/carry [5]), .IN4(n13505), .Q(n11064) );
  AO22X1 U4141 ( .IN1(\fadd_0_0_0_0_4/fracrcloseymx [5]), .IN2(n14110), .IN3(
        \fadd_0_0_0_0_4/fracrclosexmy [5]), .IN4(n14647), .Q(
        \fadd_0_0_0_0_4/fracrclose1 [5]) );
  AO22X1 U4142 ( .IN1(\fadd_0_0_0_0_4/fracrcloseymx [4]), .IN2(n14110), .IN3(
        \fadd_0_0_0_0_4/fracrclosexmy [4]), .IN4(n14647), .Q(
        \fadd_0_0_0_0_4/fracrclose1 [4]) );
  AO22X1 U4143 ( .IN1(\fadd_0_0_0_0_4/fracrcloseymx [3]), .IN2(n14110), .IN3(
        \fadd_0_0_0_0_4/fracrclosexmy [3]), .IN4(n14647), .Q(
        \fadd_0_0_0_0_4/fracrclose1 [3]) );
  AO22X1 U4144 ( .IN1(\fadd_0_0_0_0_4/fracrcloseymx [2]), .IN2(n14110), .IN3(
        \fadd_0_0_0_0_4/fracrclosexmy [2]), .IN4(n14647), .Q(
        \fadd_0_0_0_0_4/fracrclose1 [2]) );
  AO22X1 U4145 ( .IN1(\fadd_0_0_0_0_4/fracrcloseymx [1]), .IN2(n14110), .IN3(
        \fadd_0_0_0_0_4/fracrclosexmy [1]), .IN4(n14647), .Q(
        \fadd_0_0_0_0_4/fracrclose1 [1]) );
  AO22X1 U4146 ( .IN1(\fadd_0_0_0_0_4/fracrcloseymx [0]), .IN2(n14110), .IN3(
        \fadd_0_0_0_0_4/fracrcloseymx [0]), .IN4(n14647), .Q(
        \fadd_0_0_0_0_4/fracrclose1 [0]) );
  NOR3X0 U4150 ( .IN1(n14956), .IN2(n11531), .IN3(n11000), .QN(
        \fadd_0_0_0_0_4/cinaddfar ) );
  AND2X1 U4151 ( .IN1(\fadd_0_0_0_0_4/rightshiftercomponent/level1_d2[0] ), 
        .IN2(\fadd_0_0_0_0_4/rightshiftercomponent/ps_d2[0] ), .Q(n11000) );
  NOR3X0 U4153 ( .IN1(n14931), .IN2(n11529), .IN3(n10413), .QN(
        \fadd_0_0_0_0_3/zerofromclose ) );
  NAND3X0 U4155 ( .IN1(n13681), .IN2(n13489), .IN3(n11074), .QN(n11071) );
  NAND3X0 U4156 ( .IN1(n11075), .IN2(n11076), .IN3(n12841), .QN(n11070) );
  AO222X1 U4161 ( .IN1(\fadd_0_0_0_0_3/fracresultfar0 [1]), .IN2(n14743), 
        .IN3(\fadd_0_0_0_0_3/fracresultfar0 [2]), .IN4(n11080), .IN5(
        \fadd_0_0_0_0_3/fracresultfar0 [0]), .IN6(n14227), .Q(n11075) );
  AO22X1 U4162 ( .IN1(n11084), .IN2(
        \fadd_0_0_0_0_3/rightshiftercomponent/ps_d1 [1]), .IN3(n11085), .IN4(
        \fadd_0_0_0_0_3/rightshiftercomponent/ps_d1 [2]), .Q(
        \fadd_0_0_0_0_3/rightshiftercomponent/n389_o ) );
  AO22X1 U4165 ( .IN1(n13650), .IN2(\fadd_0_0_0_0_3/exponentresultclose_d1 [5]), .IN3(\fadd_0_0_0_0_3/exponentresultfar1 [5]), .IN4(n12841), .Q(
        \fadd_0_0_0_0_3/resultbeforeround [9]) );
  AO22X1 U4166 ( .IN1(n13650), .IN2(\fadd_0_0_0_0_3/exponentresultclose_d1 [4]), .IN3(\fadd_0_0_0_0_3/exponentresultfar1 [4]), .IN4(n12841), .Q(
        \fadd_0_0_0_0_3/resultbeforeround [8]) );
  AO22X1 U4167 ( .IN1(n13650), .IN2(\fadd_0_0_0_0_3/exponentresultclose_d1 [3]), .IN3(\fadd_0_0_0_0_3/exponentresultfar1 [3]), .IN4(n12841), .Q(
        \fadd_0_0_0_0_3/resultbeforeround [7]) );
  AO22X1 U4168 ( .IN1(n13650), .IN2(\fadd_0_0_0_0_3/exponentresultclose_d1 [2]), .IN3(\fadd_0_0_0_0_3/exponentresultfar1 [2]), .IN4(n12841), .Q(
        \fadd_0_0_0_0_3/resultbeforeround [6]) );
  AO22X1 U4169 ( .IN1(n13650), .IN2(\fadd_0_0_0_0_3/exponentresultclose_d1 [1]), .IN3(\fadd_0_0_0_0_3/exponentresultfar1 [1]), .IN4(n12841), .Q(
        \fadd_0_0_0_0_3/resultbeforeround [5]) );
  AO22X1 U4170 ( .IN1(n13650), .IN2(\fadd_0_0_0_0_3/exponentresultclose_d1 [0]), .IN3(\fadd_0_0_0_0_3/exponentresultfar1 [0]), .IN4(n12841), .Q(
        \fadd_0_0_0_0_3/resultbeforeround [4]) );
  AO222X1 U4171 ( .IN1(n11074), .IN2(\fadd_0_0_0_0_3/norm/level1_d1[4] ), 
        .IN3(n11087), .IN4(n13702), .IN5(n12841), .IN6(n11089), .Q(
        \fadd_0_0_0_0_3/resultbeforeround [3]) );
  AO222X1 U4172 ( .IN1(\fadd_0_0_0_0_3/fracresultfar0 [5]), .IN2(n14743), 
        .IN3(n11080), .IN4(\fadd_0_0_0_0_3/fracresultfar0 [6]), .IN5(
        \fadd_0_0_0_0_3/fracresultfar0 [4]), .IN6(n14227), .Q(n11089) );
  AO222X1 U4173 ( .IN1(n11074), .IN2(n13702), .IN3(n11087), .IN4(n13566), 
        .IN5(n12841), .IN6(n11091), .Q(\fadd_0_0_0_0_3/resultbeforeround [2])
         );
  AO222X1 U4174 ( .IN1(\fadd_0_0_0_0_3/fracresultfar0 [4]), .IN2(n14743), 
        .IN3(\fadd_0_0_0_0_3/fracresultfar0 [5]), .IN4(n11080), .IN5(n14227), 
        .IN6(\fadd_0_0_0_0_3/fracresultfar0 [3]), .Q(n11091) );
  AO222X1 U4176 ( .IN1(n11074), .IN2(n13566), .IN3(n11087), .IN4(n13489), 
        .IN5(n12841), .IN6(n11092), .Q(\fadd_0_0_0_0_3/resultbeforeround [1])
         );
  AO222X1 U4177 ( .IN1(\fadd_0_0_0_0_3/fracresultfar0 [3]), .IN2(n14743), 
        .IN3(\fadd_0_0_0_0_3/fracresultfar0 [4]), .IN4(n11080), .IN5(n14227), 
        .IN6(\fadd_0_0_0_0_3/fracresultfar0 [2]), .Q(n11092) );
  AO22X1 U4179 ( .IN1(n13650), .IN2(\fadd_0_0_0_0_3/exponentresultclose_d1 [6]), .IN3(\fadd_0_0_0_0_3/exponentresultfar1 [6]), .IN4(n12841), .Q(
        \fadd_0_0_0_0_3/resultbeforeround [10]) );
  AO222X1 U4180 ( .IN1(n11074), .IN2(n13489), .IN3(n11087), .IN4(n13681), 
        .IN5(n12841), .IN6(n11082), .Q(\fadd_0_0_0_0_3/resultbeforeround [0])
         );
  AO222X1 U4181 ( .IN1(\fadd_0_0_0_0_3/fracresultfar0 [2]), .IN2(n14743), 
        .IN3(\fadd_0_0_0_0_3/fracresultfar0 [3]), .IN4(n11080), .IN5(
        \fadd_0_0_0_0_3/fracresultfar0 [1]), .IN6(n14227), .Q(n11082) );
  AND2X1 U4188 ( .IN1(n12855), .IN2(n13650), .Q(n11074) );
  OA221X1 U4190 ( .IN1(n11093), .IN2(n11094), .IN3(n11095), .IN4(n11096), 
        .IN5(n11097), .Q(\fadd_0_0_0_0_3/ressign ) );
  XOR2X1 U4191 ( .IN1(n11098), .IN2(n11099), .Q(n11097) );
  OR3X1 U4192 ( .IN1(\fadd_0_0_0_0_3/fracrcloseymx [0]), .IN2(
        \fadd_0_0_0_0_3/fracrcloseymx [1]), .IN3(n11098), .Q(n11096) );
  OR4X1 U4195 ( .IN1(\fadd_0_0_0_0_3/fracrcloseymx [2]), .IN2(
        \fadd_0_0_0_0_3/fracrcloseymx [3]), .IN3(
        \fadd_0_0_0_0_3/fracrcloseymx [4]), .IN4(
        \fadd_0_0_0_0_3/fracrcloseymx [5]), .Q(n11095) );
  OR4X1 U4196 ( .IN1(n11100), .IN2(\fadd_0_0_0_0_3/fracrcloseymx [0]), .IN3(
        \fadd_0_0_0_0_3/fracrclosexmy [1]), .IN4(
        \fadd_0_0_0_0_3/fracrclosexmy [2]), .Q(n11094) );
  AO21X1 U4197 ( .IN1(n11101), .IN2(n11102), .IN3(n14731), .Q(n11100) );
  NAND4X0 U4198 ( .IN1(n11104), .IN2(n11105), .IN3(n14739), .IN4(n14738), .QN(
        n11102) );
  NAND4X0 U4199 ( .IN1(n11108), .IN2(n14306), .IN3(n14741), .IN4(n14740), .QN(
        n11101) );
  AO21X1 U4201 ( .IN1(\fadd_0_0_0_0_3/sub_784/B[1] ), .IN2(n14051), .IN3(
        n11113), .Q(\fadd_0_0_0_0_3/norm/level1 [4]) );
  OAI22X1 U4203 ( .IN1(n14931), .IN2(n11520), .IN3(n11114), .IN4(n11897), .QN(
        \fadd_0_0_0_0_3/norm/level1 [3]) );
  OAI22X1 U4204 ( .IN1(n14931), .IN2(n11519), .IN3(n11114), .IN4(n11898), .QN(
        \fadd_0_0_0_0_3/norm/level1 [2]) );
  NOR3X0 U4209 ( .IN1(n13545), .IN2(n8644), .IN3(n11113), .QN(
        \fadd_0_0_0_0_3/sub_784/B[1] ) );
  OAI21X1 U4210 ( .IN1(n10413), .IN2(n11519), .IN3(n11896), .QN(n11113) );
  NAND4X0 U4213 ( .IN1(n11895), .IN2(n11896), .IN3(n11897), .IN4(n11898), .QN(
        n10413) );
  AO22X1 U4214 ( .IN1(n14306), .IN2(n13510), .IN3(n11105), .IN4(n13623), .Q(
        \fadd_0_0_0_0_3/newy_11 ) );
  AO22X1 U4215 ( .IN1(n14306), .IN2(n13474), .IN3(n11105), .IN4(n13890), .Q(
        \fadd_0_0_0_0_3/newy_10 ) );
  AO22X1 U4216 ( .IN1(n14306), .IN2(n5770), .IN3(n11105), .IN4(n5782), .Q(
        \fadd_0_0_0_0_3/newx [8]) );
  AO22X1 U4219 ( .IN1(n14306), .IN2(n5769), .IN3(n11105), .IN4(n5781), .Q(
        \fadd_0_0_0_0_3/newx [7]) );
  AO22X1 U4222 ( .IN1(n14306), .IN2(n5768), .IN3(n11105), .IN4(n5780), .Q(
        \fadd_0_0_0_0_3/newx [6]) );
  AO22X1 U4225 ( .IN1(n14306), .IN2(n5767), .IN3(n11105), .IN4(n5779), .Q(
        \fadd_0_0_0_0_3/newx [5]) );
  AO22X1 U4228 ( .IN1(n14306), .IN2(n5766), .IN3(n11105), .IN4(n5778), .Q(
        \fadd_0_0_0_0_3/newx [4]) );
  AO22X1 U4231 ( .IN1(n14306), .IN2(n13709), .IN3(n11105), .IN4(n13571), .Q(
        \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ) );
  AO22X1 U4234 ( .IN1(n14306), .IN2(n13687), .IN3(n11105), .IN4(n13554), .Q(
        \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ) );
  AO22X1 U4237 ( .IN1(n14306), .IN2(n13666), .IN3(n11105), .IN4(n13529), .Q(
        \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ) );
  AO22X1 U4241 ( .IN1(n14306), .IN2(n13890), .IN3(n11105), .IN4(n13474), .Q(
        \fadd_0_0_0_0_3/newx [10]) );
  AO22X1 U4243 ( .IN1(n14306), .IN2(n13638), .IN3(n11105), .IN4(n13518), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ) );
  XOR2X1 U4246 ( .IN1(n11115), .IN2(n14731), .Q(
        \fadd_0_0_0_0_3/fracyfarxorop [6]) );
  XOR2X1 U4248 ( .IN1(n11118), .IN2(n12722), .Q(
        \fadd_0_0_0_0_3/fracyfarxorop [5]) );
  OA21X1 U4249 ( .IN1(n12719), .IN2(n14733), .IN3(n14728), .Q(n11118) );
  XOR2X1 U4251 ( .IN1(n11121), .IN2(n12722), .Q(
        \fadd_0_0_0_0_3/fracyfarxorop [4]) );
  OA22X1 U4252 ( .IN1(n14730), .IN2(n11122), .IN3(n12719), .IN4(n11123), .Q(
        n11121) );
  AO22X1 U4254 ( .IN1(n11125), .IN2(n14730), .IN3(n11126), .IN4(n12719), .Q(
        \fadd_0_0_0_0_3/fracyfarxorop [3]) );
  XOR2X1 U4255 ( .IN1(n11123), .IN2(n12722), .Q(n11126) );
  AO21X1 U4256 ( .IN1(n14734), .IN2(n11128), .IN3(n14727), .Q(n11123) );
  AO22X1 U4257 ( .IN1(n11130), .IN2(n14730), .IN3(n11125), .IN4(n12719), .Q(
        \fadd_0_0_0_0_3/fracyfarxorop [2]) );
  XOR2X1 U4258 ( .IN1(n14731), .IN2(n11131), .Q(n11125) );
  OA22X1 U4259 ( .IN1(n11124), .IN2(n11132), .IN3(n11133), .IN4(n11120), .Q(
        n11131) );
  AO22X1 U4261 ( .IN1(n11135), .IN2(n14730), .IN3(n11130), .IN4(n12719), .Q(
        \fadd_0_0_0_0_3/fracyfarxorop [1]) );
  XOR2X1 U4262 ( .IN1(n14731), .IN2(n11136), .Q(n11130) );
  OA22X1 U4263 ( .IN1(n11137), .IN2(n11132), .IN3(n14729), .IN4(n11138), .Q(
        n11136) );
  AO22X1 U4265 ( .IN1(n11135), .IN2(n12719), .IN3(n11139), .IN4(n14730), .Q(
        \fadd_0_0_0_0_3/fracyfarxorop [0]) );
  XOR2X1 U4267 ( .IN1(n12720), .IN2(n12722), .Q(n11139) );
  OA22X1 U4268 ( .IN1(n14729), .IN2(n12721), .IN3(n14736), .IN4(n14726), .Q(
        n12720) );
  XOR2X1 U4272 ( .IN1(n14731), .IN2(n11141), .Q(n11135) );
  AOI22X1 U4273 ( .IN1(n14735), .IN2(n14727), .IN3(n11134), .IN4(
        \fadd_0_0_0_0_3/rightshiftercomponent/level2[1] ), .QN(n11141) );
  OA221X1 U4277 ( .IN1(n14738), .IN2(n14306), .IN3(n14740), .IN4(n11105), 
        .IN5(n11140), .Q(n11128) );
  OA221X1 U4281 ( .IN1(n14739), .IN2(n14306), .IN3(n14741), .IN4(n11105), 
        .IN5(n11140), .Q(n11134) );
  OA22X1 U4282 ( .IN1(n14306), .IN2(n11104), .IN3(n11108), .IN4(n11105), .Q(
        n11140) );
  XOR2X1 U4288 ( .IN1(n14732), .IN2(\fadd_0_0_0_0_3/newy_9 ), .Q(n12722) );
  AO22X1 U4289 ( .IN1(n14306), .IN2(n13580), .IN3(n11105), .IN4(n13718), .Q(
        \fadd_0_0_0_0_3/newy_9 ) );
  OA22X1 U4293 ( .IN1(n11105), .IN2(n11686), .IN3(n14306), .IN4(n11697), .Q(
        n11099) );
  AO22X1 U4295 ( .IN1(n14737), .IN2(n14734), .IN3(n14733), .IN4(n11142), .Q(
        \fadd_0_0_0_0_3/fracyclose1 [3]) );
  OA22X1 U4297 ( .IN1(n11105), .IN2(n11691), .IN3(n14306), .IN4(n11680), .Q(
        n11124) );
  AO22X1 U4298 ( .IN1(n14737), .IN2(n14735), .IN3(n14734), .IN4(n11142), .Q(
        \fadd_0_0_0_0_3/fracyclose1 [2]) );
  OA22X1 U4300 ( .IN1(n11105), .IN2(n11690), .IN3(n14306), .IN4(n11679), .Q(
        n11137) );
  AO22X1 U4301 ( .IN1(n14735), .IN2(n11142), .IN3(n14737), .IN4(n14736), .Q(
        \fadd_0_0_0_0_3/fracyclose1 [1]) );
  OA22X1 U4304 ( .IN1(n11105), .IN2(n11689), .IN3(n14306), .IN4(n11678), .Q(
        n11133) );
  OA22X1 U4306 ( .IN1(n11105), .IN2(n11688), .IN3(n14306), .IN4(n11677), .Q(
        n11143) );
  AO22X1 U4308 ( .IN1(\fadd_0_0_0_0_3/exponentdifferenceyx [0]), .IN2(n14306), 
        .IN3(\fadd_0_0_0_0_3/exponentdifferencexy [0]), .IN4(n11105), .Q(
        n11142) );
  OA22X1 U4311 ( .IN1(n11687), .IN2(n11146), .IN3(
        \fadd_0_0_0_0_3/sub_707/carry [5]), .IN4(n13474), .Q(n11145) );
  AO22X1 U4318 ( .IN1(\fadd_0_0_0_0_3/fracrcloseymx [5]), .IN2(n14117), .IN3(
        \fadd_0_0_0_0_3/fracrclosexmy [5]), .IN4(n14642), .Q(
        \fadd_0_0_0_0_3/fracrclose1 [5]) );
  AO22X1 U4319 ( .IN1(\fadd_0_0_0_0_3/fracrcloseymx [4]), .IN2(n14117), .IN3(
        \fadd_0_0_0_0_3/fracrclosexmy [4]), .IN4(n14642), .Q(
        \fadd_0_0_0_0_3/fracrclose1 [4]) );
  AO22X1 U4320 ( .IN1(\fadd_0_0_0_0_3/fracrcloseymx [3]), .IN2(n14117), .IN3(
        \fadd_0_0_0_0_3/fracrclosexmy [3]), .IN4(n14642), .Q(
        \fadd_0_0_0_0_3/fracrclose1 [3]) );
  AO22X1 U4321 ( .IN1(\fadd_0_0_0_0_3/fracrcloseymx [2]), .IN2(n14117), .IN3(
        \fadd_0_0_0_0_3/fracrclosexmy [2]), .IN4(n14642), .Q(
        \fadd_0_0_0_0_3/fracrclose1 [2]) );
  AO22X1 U4322 ( .IN1(\fadd_0_0_0_0_3/fracrcloseymx [1]), .IN2(n14117), .IN3(
        \fadd_0_0_0_0_3/fracrclosexmy [1]), .IN4(n14642), .Q(
        \fadd_0_0_0_0_3/fracrclose1 [1]) );
  AO22X1 U4323 ( .IN1(\fadd_0_0_0_0_3/fracrcloseymx [0]), .IN2(n14117), .IN3(
        \fadd_0_0_0_0_3/fracrcloseymx [0]), .IN4(n14642), .Q(
        \fadd_0_0_0_0_3/fracrclose1 [0]) );
  NOR3X0 U4327 ( .IN1(n14947), .IN2(n11518), .IN3(n11081), .QN(
        \fadd_0_0_0_0_3/cinaddfar ) );
  AND2X1 U4328 ( .IN1(\fadd_0_0_0_0_3/rightshiftercomponent/level1_d2[0] ), 
        .IN2(\fadd_0_0_0_0_3/rightshiftercomponent/ps_d2[0] ), .Q(n11081) );
  NOR3X0 U4330 ( .IN1(n14930), .IN2(n11516), .IN3(n10412), .QN(
        \fadd_0_0_0_0_2/zerofromclose ) );
  NAND3X0 U4332 ( .IN1(n13675), .IN2(n13484), .IN3(n11155), .QN(n11152) );
  NAND3X0 U4333 ( .IN1(n11156), .IN2(n11157), .IN3(n12840), .QN(n11151) );
  AO222X1 U4338 ( .IN1(\fadd_0_0_0_0_2/fracresultfar0 [1]), .IN2(n14722), 
        .IN3(\fadd_0_0_0_0_2/fracresultfar0 [2]), .IN4(n11161), .IN5(
        \fadd_0_0_0_0_2/fracresultfar0 [0]), .IN6(n14226), .Q(n11156) );
  AO22X1 U4339 ( .IN1(n11165), .IN2(
        \fadd_0_0_0_0_2/rightshiftercomponent/ps_d1 [1]), .IN3(n11166), .IN4(
        \fadd_0_0_0_0_2/rightshiftercomponent/ps_d1 [2]), .Q(
        \fadd_0_0_0_0_2/rightshiftercomponent/n389_o ) );
  AO22X1 U4342 ( .IN1(n13645), .IN2(\fadd_0_0_0_0_2/exponentresultclose_d1 [5]), .IN3(\fadd_0_0_0_0_2/exponentresultfar1 [5]), .IN4(n12840), .Q(
        \fadd_0_0_0_0_2/resultbeforeround [9]) );
  AO22X1 U4343 ( .IN1(n13645), .IN2(\fadd_0_0_0_0_2/exponentresultclose_d1 [4]), .IN3(\fadd_0_0_0_0_2/exponentresultfar1 [4]), .IN4(n12840), .Q(
        \fadd_0_0_0_0_2/resultbeforeround [8]) );
  AO22X1 U4344 ( .IN1(n13645), .IN2(\fadd_0_0_0_0_2/exponentresultclose_d1 [3]), .IN3(\fadd_0_0_0_0_2/exponentresultfar1 [3]), .IN4(n12840), .Q(
        \fadd_0_0_0_0_2/resultbeforeround [7]) );
  AO22X1 U4345 ( .IN1(n13645), .IN2(\fadd_0_0_0_0_2/exponentresultclose_d1 [2]), .IN3(\fadd_0_0_0_0_2/exponentresultfar1 [2]), .IN4(n12840), .Q(
        \fadd_0_0_0_0_2/resultbeforeround [6]) );
  AO22X1 U4346 ( .IN1(n13645), .IN2(\fadd_0_0_0_0_2/exponentresultclose_d1 [1]), .IN3(\fadd_0_0_0_0_2/exponentresultfar1 [1]), .IN4(n12840), .Q(
        \fadd_0_0_0_0_2/resultbeforeround [5]) );
  AO22X1 U4347 ( .IN1(n13645), .IN2(\fadd_0_0_0_0_2/exponentresultclose_d1 [0]), .IN3(\fadd_0_0_0_0_2/exponentresultfar1 [0]), .IN4(n12840), .Q(
        \fadd_0_0_0_0_2/resultbeforeround [4]) );
  AO222X1 U4348 ( .IN1(n11155), .IN2(\fadd_0_0_0_0_2/norm/level1_d1[4] ), 
        .IN3(n11168), .IN4(n13694), .IN5(n12840), .IN6(n11170), .Q(
        \fadd_0_0_0_0_2/resultbeforeround [3]) );
  AO222X1 U4349 ( .IN1(\fadd_0_0_0_0_2/fracresultfar0 [5]), .IN2(n14722), 
        .IN3(n11161), .IN4(\fadd_0_0_0_0_2/fracresultfar0 [6]), .IN5(
        \fadd_0_0_0_0_2/fracresultfar0 [4]), .IN6(n14226), .Q(n11170) );
  AO222X1 U4350 ( .IN1(n11155), .IN2(n13694), .IN3(n11168), .IN4(n13552), 
        .IN5(n12840), .IN6(n11172), .Q(\fadd_0_0_0_0_2/resultbeforeround [2])
         );
  AO222X1 U4351 ( .IN1(\fadd_0_0_0_0_2/fracresultfar0 [4]), .IN2(n14722), 
        .IN3(\fadd_0_0_0_0_2/fracresultfar0 [5]), .IN4(n11161), .IN5(n14226), 
        .IN6(\fadd_0_0_0_0_2/fracresultfar0 [3]), .Q(n11172) );
  AO222X1 U4353 ( .IN1(n11155), .IN2(n13552), .IN3(n11168), .IN4(n13484), 
        .IN5(n12840), .IN6(n11173), .Q(\fadd_0_0_0_0_2/resultbeforeround [1])
         );
  AO222X1 U4354 ( .IN1(\fadd_0_0_0_0_2/fracresultfar0 [3]), .IN2(n14722), 
        .IN3(\fadd_0_0_0_0_2/fracresultfar0 [4]), .IN4(n11161), .IN5(n14226), 
        .IN6(\fadd_0_0_0_0_2/fracresultfar0 [2]), .Q(n11173) );
  AO22X1 U4356 ( .IN1(n13645), .IN2(\fadd_0_0_0_0_2/exponentresultclose_d1 [6]), .IN3(\fadd_0_0_0_0_2/exponentresultfar1 [6]), .IN4(n12840), .Q(
        \fadd_0_0_0_0_2/resultbeforeround [10]) );
  AO222X1 U4357 ( .IN1(n11155), .IN2(n13484), .IN3(n11168), .IN4(n13675), 
        .IN5(n12840), .IN6(n11163), .Q(\fadd_0_0_0_0_2/resultbeforeround [0])
         );
  AO222X1 U4358 ( .IN1(\fadd_0_0_0_0_2/fracresultfar0 [2]), .IN2(n14722), 
        .IN3(\fadd_0_0_0_0_2/fracresultfar0 [3]), .IN4(n11161), .IN5(
        \fadd_0_0_0_0_2/fracresultfar0 [1]), .IN6(n14226), .Q(n11163) );
  AND2X1 U4365 ( .IN1(n12853), .IN2(n13645), .Q(n11155) );
  OA221X1 U4367 ( .IN1(n11174), .IN2(n11175), .IN3(n11176), .IN4(n11177), 
        .IN5(n11178), .Q(\fadd_0_0_0_0_2/ressign ) );
  OR4X1 U4372 ( .IN1(\fadd_0_0_0_0_2/fracrcloseymx [2]), .IN2(
        \fadd_0_0_0_0_2/fracrcloseymx [3]), .IN3(
        \fadd_0_0_0_0_2/fracrcloseymx [4]), .IN4(
        \fadd_0_0_0_0_2/fracrcloseymx [5]), .Q(n11176) );
  OR4X1 U4373 ( .IN1(n11181), .IN2(\fadd_0_0_0_0_2/fracrcloseymx [0]), .IN3(
        \fadd_0_0_0_0_2/fracrclosexmy [1]), .IN4(
        \fadd_0_0_0_0_2/fracrclosexmy [2]), .Q(n11175) );
  AO21X1 U4374 ( .IN1(n11182), .IN2(n11183), .IN3(n14699), .Q(n11181) );
  NAND4X0 U4375 ( .IN1(n11185), .IN2(n11186), .IN3(n14707), .IN4(n14706), .QN(
        n11183) );
  NAND4X0 U4376 ( .IN1(n11189), .IN2(n14305), .IN3(n14709), .IN4(n14708), .QN(
        n11182) );
  AO21X1 U4378 ( .IN1(\fadd_0_0_0_0_2/sub_784/B[1] ), .IN2(n14050), .IN3(
        n11194), .Q(\fadd_0_0_0_0_2/norm/level1 [4]) );
  OAI22X1 U4380 ( .IN1(n14930), .IN2(n11507), .IN3(n11195), .IN4(n11893), .QN(
        \fadd_0_0_0_0_2/norm/level1 [3]) );
  OAI22X1 U4381 ( .IN1(n14930), .IN2(n11506), .IN3(n11195), .IN4(n11894), .QN(
        \fadd_0_0_0_0_2/norm/level1 [2]) );
  NOR3X0 U4386 ( .IN1(n13546), .IN2(n8640), .IN3(n11194), .QN(
        \fadd_0_0_0_0_2/sub_784/B[1] ) );
  OAI21X1 U4387 ( .IN1(n10412), .IN2(n11506), .IN3(n11892), .QN(n11194) );
  NAND4X0 U4390 ( .IN1(n11891), .IN2(n11892), .IN3(n11893), .IN4(n11894), .QN(
        n10412) );
  AO22X1 U4391 ( .IN1(n14305), .IN2(n13507), .IN3(n11186), .IN4(n13470), .Q(
        \fadd_0_0_0_0_2/newy_11 ) );
  AO22X1 U4392 ( .IN1(n14305), .IN2(n13472), .IN3(n11186), .IN4(n13589), .Q(
        \fadd_0_0_0_0_2/newy_10 ) );
  AO22X1 U4393 ( .IN1(n14305), .IN2(n5842), .IN3(n11186), .IN4(n5854), .Q(
        \fadd_0_0_0_0_2/newx [8]) );
  AO22X1 U4396 ( .IN1(n14305), .IN2(n5841), .IN3(n11186), .IN4(n5853), .Q(
        \fadd_0_0_0_0_2/newx [7]) );
  AO22X1 U4399 ( .IN1(n14305), .IN2(n5840), .IN3(n11186), .IN4(n5852), .Q(
        \fadd_0_0_0_0_2/newx [6]) );
  AO22X1 U4402 ( .IN1(n14305), .IN2(n5839), .IN3(n11186), .IN4(n5851), .Q(
        \fadd_0_0_0_0_2/newx [5]) );
  AO22X1 U4405 ( .IN1(n14305), .IN2(n5838), .IN3(n11186), .IN4(n5850), .Q(
        \fadd_0_0_0_0_2/newx [4]) );
  AO22X1 U4408 ( .IN1(n14305), .IN2(n13577), .IN3(n11186), .IN4(n13495), .Q(
        \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ) );
  AO22X1 U4411 ( .IN1(n14305), .IN2(n13560), .IN3(n11186), .IN4(n13493), .Q(
        \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ) );
  AO22X1 U4414 ( .IN1(n14305), .IN2(n13535), .IN3(n11186), .IN4(n13480), .Q(
        \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ) );
  AO22X1 U4418 ( .IN1(n14305), .IN2(n13589), .IN3(n11186), .IN4(n13472), .Q(
        \fadd_0_0_0_0_2/newx [10]) );
  AO22X1 U4420 ( .IN1(n14305), .IN2(n13524), .IN3(n11186), .IN4(n13478), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ) );
  XOR2X1 U4423 ( .IN1(n11196), .IN2(n14699), .Q(
        \fadd_0_0_0_0_2/fracyfarxorop [6]) );
  XOR2X1 U4425 ( .IN1(n11199), .IN2(n12714), .Q(
        \fadd_0_0_0_0_2/fracyfarxorop [5]) );
  OA21X1 U4426 ( .IN1(n12711), .IN2(n14701), .IN3(n14696), .Q(n11199) );
  XOR2X1 U4428 ( .IN1(n11202), .IN2(n12714), .Q(
        \fadd_0_0_0_0_2/fracyfarxorop [4]) );
  OA22X1 U4429 ( .IN1(n14698), .IN2(n11203), .IN3(n12711), .IN4(n11204), .Q(
        n11202) );
  AO22X1 U4431 ( .IN1(n11206), .IN2(n14698), .IN3(n11207), .IN4(n12711), .Q(
        \fadd_0_0_0_0_2/fracyfarxorop [3]) );
  XOR2X1 U4432 ( .IN1(n11204), .IN2(n12714), .Q(n11207) );
  AO21X1 U4433 ( .IN1(n14702), .IN2(n11209), .IN3(n14695), .Q(n11204) );
  AO22X1 U4434 ( .IN1(n11211), .IN2(n14698), .IN3(n11206), .IN4(n12711), .Q(
        \fadd_0_0_0_0_2/fracyfarxorop [2]) );
  XOR2X1 U4435 ( .IN1(n14699), .IN2(n11212), .Q(n11206) );
  OA22X1 U4436 ( .IN1(n11205), .IN2(n11213), .IN3(n11214), .IN4(n11201), .Q(
        n11212) );
  AO22X1 U4438 ( .IN1(n11216), .IN2(n14698), .IN3(n11211), .IN4(n12711), .Q(
        \fadd_0_0_0_0_2/fracyfarxorop [1]) );
  XOR2X1 U4439 ( .IN1(n14699), .IN2(n11217), .Q(n11211) );
  OA22X1 U4440 ( .IN1(n11218), .IN2(n11213), .IN3(n14697), .IN4(n11219), .Q(
        n11217) );
  AO22X1 U4442 ( .IN1(n11216), .IN2(n12711), .IN3(n11220), .IN4(n14698), .Q(
        \fadd_0_0_0_0_2/fracyfarxorop [0]) );
  XOR2X1 U4444 ( .IN1(n12712), .IN2(n12714), .Q(n11220) );
  OA22X1 U4445 ( .IN1(n14697), .IN2(n12713), .IN3(n14704), .IN4(n14694), .Q(
        n12712) );
  XOR2X1 U4449 ( .IN1(n14699), .IN2(n11222), .Q(n11216) );
  AOI22X1 U4450 ( .IN1(n14703), .IN2(n14695), .IN3(n11215), .IN4(
        \fadd_0_0_0_0_2/rightshiftercomponent/level2[1] ), .QN(n11222) );
  OA221X1 U4454 ( .IN1(n14706), .IN2(n14305), .IN3(n14708), .IN4(n11186), 
        .IN5(n11221), .Q(n11209) );
  OA221X1 U4458 ( .IN1(n14707), .IN2(n14305), .IN3(n14709), .IN4(n11186), 
        .IN5(n11221), .Q(n11215) );
  OA22X1 U4459 ( .IN1(n14305), .IN2(n11185), .IN3(n11189), .IN4(n11186), .Q(
        n11221) );
  XOR2X1 U4465 ( .IN1(n14700), .IN2(\fadd_0_0_0_0_2/newy_9 ), .Q(n12714) );
  OAI22X1 U4466 ( .IN1(n11186), .IN2(n11718), .IN3(n14305), .IN4(n11707), .QN(
        \fadd_0_0_0_0_2/newy_9 ) );
  OA22X1 U4468 ( .IN1(n11186), .IN2(n11707), .IN3(n14305), .IN4(n11718), .Q(
        n11180) );
  AO22X1 U4470 ( .IN1(n14705), .IN2(n14702), .IN3(n14701), .IN4(n11223), .Q(
        \fadd_0_0_0_0_2/fracyclose1 [3]) );
  OA22X1 U4472 ( .IN1(n11186), .IN2(n11712), .IN3(n14305), .IN4(n11701), .Q(
        n11205) );
  AO22X1 U4473 ( .IN1(n14705), .IN2(n14703), .IN3(n14702), .IN4(n11223), .Q(
        \fadd_0_0_0_0_2/fracyclose1 [2]) );
  OA22X1 U4475 ( .IN1(n11186), .IN2(n11711), .IN3(n14305), .IN4(n11700), .Q(
        n11218) );
  AO22X1 U4476 ( .IN1(n14703), .IN2(n11223), .IN3(n14705), .IN4(n14704), .Q(
        \fadd_0_0_0_0_2/fracyclose1 [1]) );
  OA22X1 U4479 ( .IN1(n11186), .IN2(n11710), .IN3(n14305), .IN4(n11699), .Q(
        n11214) );
  OA22X1 U4481 ( .IN1(n11186), .IN2(n11709), .IN3(n14305), .IN4(n11698), .Q(
        n11224) );
  AO22X1 U4483 ( .IN1(\fadd_0_0_0_0_2/exponentdifferenceyx [0]), .IN2(n14305), 
        .IN3(\fadd_0_0_0_0_2/exponentdifferencexy [0]), .IN4(n11186), .Q(
        n11223) );
  OA22X1 U4486 ( .IN1(n11708), .IN2(n11227), .IN3(
        \fadd_0_0_0_0_2/sub_707/carry [5]), .IN4(n13472), .Q(n11226) );
  AO22X1 U4493 ( .IN1(\fadd_0_0_0_0_2/fracrcloseymx [5]), .IN2(n14112), .IN3(
        \fadd_0_0_0_0_2/fracrclosexmy [5]), .IN4(n14643), .Q(
        \fadd_0_0_0_0_2/fracrclose1 [5]) );
  AO22X1 U4494 ( .IN1(\fadd_0_0_0_0_2/fracrcloseymx [4]), .IN2(n14112), .IN3(
        \fadd_0_0_0_0_2/fracrclosexmy [4]), .IN4(n14643), .Q(
        \fadd_0_0_0_0_2/fracrclose1 [4]) );
  AO22X1 U4495 ( .IN1(\fadd_0_0_0_0_2/fracrcloseymx [3]), .IN2(n14112), .IN3(
        \fadd_0_0_0_0_2/fracrclosexmy [3]), .IN4(n14643), .Q(
        \fadd_0_0_0_0_2/fracrclose1 [3]) );
  AO22X1 U4496 ( .IN1(\fadd_0_0_0_0_2/fracrcloseymx [2]), .IN2(n14112), .IN3(
        \fadd_0_0_0_0_2/fracrclosexmy [2]), .IN4(n14643), .Q(
        \fadd_0_0_0_0_2/fracrclose1 [2]) );
  AO22X1 U4497 ( .IN1(\fadd_0_0_0_0_2/fracrcloseymx [1]), .IN2(n14112), .IN3(
        \fadd_0_0_0_0_2/fracrclosexmy [1]), .IN4(n14643), .Q(
        \fadd_0_0_0_0_2/fracrclose1 [1]) );
  AO22X1 U4498 ( .IN1(\fadd_0_0_0_0_2/fracrcloseymx [0]), .IN2(n14112), .IN3(
        \fadd_0_0_0_0_2/fracrcloseymx [0]), .IN4(n14643), .Q(
        \fadd_0_0_0_0_2/fracrclose1 [0]) );
  NOR3X0 U4502 ( .IN1(n14946), .IN2(n11505), .IN3(n11162), .QN(
        \fadd_0_0_0_0_2/cinaddfar ) );
  AND2X1 U4503 ( .IN1(\fadd_0_0_0_0_2/rightshiftercomponent/level1_d2[0] ), 
        .IN2(\fadd_0_0_0_0_2/rightshiftercomponent/ps_d2[0] ), .Q(n11162) );
  AO22X1 U4505 ( .IN1(n11232), .IN2(
        \fadd_0_0_0_0_10/rightshiftercomponent/n43 ), .IN3(n11233), .IN4(
        \fadd_0_0_0_0_10/rightshiftercomponent/n44 ), .Q(
        \fadd_0_0_0_0_10/rightshiftercomponent/n11 ) );
  NAND3X0 U4509 ( .IN1(n11235), .IN2(n11236), .IN3(n11887), .QN(
        \fadd_0_0_0_0_10/norm/U5/Z_5 ) );
  OR2X1 U4510 ( .IN1(n12870), .IN2(n11889), .Q(n11235) );
  OAI21X1 U4511 ( .IN1(n12870), .IN2(n11890), .IN3(n11237), .QN(
        \fadd_0_0_0_0_10/norm/U5/Z_4 ) );
  OAI22X1 U4512 ( .IN1(n12870), .IN2(n11499), .IN3(n11238), .IN4(n11889), .QN(
        \fadd_0_0_0_0_10/norm/U5/Z_3 ) );
  OAI22X1 U4513 ( .IN1(n12870), .IN2(n11498), .IN3(n11238), .IN4(n11890), .QN(
        \fadd_0_0_0_0_10/norm/U5/Z_2 ) );
  XOR2X1 U4517 ( .IN1(n11239), .IN2(n11240), .Q(\fadd_0_0_0_0_10/n240 ) );
  XOR2X1 U4519 ( .IN1(n11243), .IN2(n14938), .Q(\fadd_0_0_0_0_10/n239 ) );
  OA21X1 U4520 ( .IN1(n14978), .IN2(n14974), .IN3(n11241), .Q(n11243) );
  XOR2X1 U4521 ( .IN1(n11245), .IN2(n14938), .Q(\fadd_0_0_0_0_10/n238 ) );
  OA22X1 U4522 ( .IN1(n11242), .IN2(n11246), .IN3(n14978), .IN4(n11247), .Q(
        n11245) );
  AO22X1 U4524 ( .IN1(n11249), .IN2(n11242), .IN3(n11250), .IN4(n14978), .Q(
        \fadd_0_0_0_0_10/n237 ) );
  XOR2X1 U4525 ( .IN1(n11247), .IN2(n14938), .Q(n11250) );
  OAI21X1 U4526 ( .IN1(n11251), .IN2(\fadd_0_0_0_0_10/U27/Z_2 ), .IN3(n11252), 
        .QN(n11247) );
  AO22X1 U4527 ( .IN1(n11253), .IN2(n11242), .IN3(n11249), .IN4(n14978), .Q(
        \fadd_0_0_0_0_10/n236 ) );
  XOR2X1 U4528 ( .IN1(n11240), .IN2(n11254), .Q(n11249) );
  OA22X1 U4529 ( .IN1(n10409), .IN2(n11252), .IN3(n11255), .IN4(n14977), .Q(
        n11254) );
  AO22X1 U4532 ( .IN1(n11256), .IN2(n11242), .IN3(n11253), .IN4(n14978), .Q(
        \fadd_0_0_0_0_10/n235 ) );
  XOR2X1 U4533 ( .IN1(n11240), .IN2(n11257), .Q(n11253) );
  OA22X1 U4534 ( .IN1(n11251), .IN2(n11252), .IN3(\fadd_0_0_0_0_10/U27/Z_1 ), 
        .IN4(n11258), .Q(n11257) );
  AO22X1 U4536 ( .IN1(n11256), .IN2(n14978), .IN3(n11259), .IN4(n11242), .Q(
        \fadd_0_0_0_0_10/n234 ) );
  XOR2X1 U4537 ( .IN1(n14938), .IN2(
        \fadd_0_0_0_0_10/rightshiftercomponent/U5/Z_0 ), .Q(n11259) );
  AO21X1 U4538 ( .IN1(n11260), .IN2(\fadd_0_0_0_0_10/U27/Z_1 ), .IN3(
        \fadd_0_0_0_0_10/rightshiftercomponent/U6/Z_0 ), .Q(
        \fadd_0_0_0_0_10/rightshiftercomponent/U5/Z_0 ) );
  XOR2X1 U4544 ( .IN1(n11240), .IN2(n11264), .Q(n11256) );
  OA22X1 U4545 ( .IN1(n11255), .IN2(n11252), .IN3(\fadd_0_0_0_0_10/U27/Z_1 ), 
        .IN4(n11234), .Q(n11264) );
  NOR3X0 U4549 ( .IN1(n12871), .IN2(n11497), .IN3(n12870), .QN(
        \fadd_0_0_0_0_10/n182 ) );
  NAND3X0 U4550 ( .IN1(n11887), .IN2(n11236), .IN3(n11237), .QN(n12870) );
  OA21X1 U4551 ( .IN1(n12871), .IN2(n11498), .IN3(n11888), .Q(n11237) );
  OR2X1 U4552 ( .IN1(n12871), .IN2(n11499), .Q(n11236) );
  NAND4X0 U4553 ( .IN1(n11887), .IN2(n11888), .IN3(n11889), .IN4(n11890), .QN(
        n12871) );
  NOR3X0 U4554 ( .IN1(n13616), .IN2(n11496), .IN3(n8883), .QN(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/CI )
         );
  AND2X1 U4555 ( .IN1(\fadd_0_0_0_0_10/rightshiftercomponent/n16 ), .IN2(
        \fadd_0_0_0_0_10/rightshiftercomponent/n41 ), .Q(n8883) );
  AOI21X1 U4557 ( .IN1(n14987), .IN2(n12067), .IN3(n14993), .QN(
        \fadd_0_0_0_0_10/add_859/carry[6] ) );
  AO22X1 U4559 ( .IN1(n13412), .IN2(n11266), .IN3(n11267), .IN4(n14988), .Q(
        n8804) );
  NAND3X0 U4562 ( .IN1(n8826), .IN2(n12028), .IN3(n12032), .QN(n11266) );
  OA21X1 U4563 ( .IN1(n14993), .IN2(n11268), .IN3(n8837), .Q(n8826) );
  AO22X1 U4572 ( .IN1(n14304), .IN2(n14983), .IN3(n11271), .IN4(n14999), .Q(
        \fadd_0_0_0_0_10/U29/Z_8 ) );
  AO22X1 U4575 ( .IN1(n14304), .IN2(n14982), .IN3(n11271), .IN4(n14998), .Q(
        \fadd_0_0_0_0_10/U29/Z_7 ) );
  AO22X1 U4578 ( .IN1(n14304), .IN2(n14981), .IN3(n11271), .IN4(n14997), .Q(
        \fadd_0_0_0_0_10/U29/Z_6 ) );
  AO22X1 U4581 ( .IN1(n14188), .IN2(n14980), .IN3(n11271), .IN4(n14996), .Q(
        \fadd_0_0_0_0_10/U29/Z_5 ) );
  AO22X1 U4584 ( .IN1(n14188), .IN2(n13885), .IN3(n11271), .IN4(n13635), .Q(
        \fadd_0_0_0_0_10/U29/Z_4 ) );
  OA22X1 U4587 ( .IN1(n13696), .IN2(n11271), .IN3(n13562), .IN4(n14304), .Q(
        \fadd_0_0_0_0_10/U29/Z_3 ) );
  OA22X1 U4590 ( .IN1(n13673), .IN2(n11271), .IN3(n13538), .IN4(n14304), .Q(
        \fadd_0_0_0_0_10/U29/Z_2 ) );
  AO22X1 U4594 ( .IN1(n14304), .IN2(n13887), .IN3(n11271), .IN4(n13469), .Q(
        \fadd_0_0_0_0_10/U29/Z_10 ) );
  OA22X1 U4595 ( .IN1(n13646), .IN2(n11271), .IN3(n13526), .IN4(n14304), .Q(
        \fadd_0_0_0_0_10/U29/Z_1 ) );
  OA22X1 U4598 ( .IN1(n13633), .IN2(n11271), .IN3(n13477), .IN4(n14304), .Q(
        \fadd_0_0_0_0_10/U29/Z_0 ) );
  AO22X1 U4601 ( .IN1(n14188), .IN2(n13500), .IN3(n11271), .IN4(n13886), .Q(
        \fadd_0_0_0_0_10/U28/Z_6 ) );
  AO22X1 U4603 ( .IN1(n14188), .IN2(n13469), .IN3(n11271), .IN4(n13887), .Q(
        \fadd_0_0_0_0_10/U28/Z_5 ) );
  OA22X1 U4608 ( .IN1(n14971), .IN2(\fadd_0_0_0_0_10/U27/DATA1_0 ), .IN3(
        n14974), .IN4(n14979), .Q(\fadd_0_0_0_0_10/U25/Z_3 ) );
  OA22X1 U4610 ( .IN1(n11271), .IN2(n11853), .IN3(n14304), .IN4(n11848), .Q(
        n10409) );
  OA22X1 U4611 ( .IN1(\fadd_0_0_0_0_10/U27/DATA1_0 ), .IN2(n14968), .IN3(
        n14971), .IN4(n14979), .Q(\fadd_0_0_0_0_10/U25/Z_2 ) );
  OA22X1 U4613 ( .IN1(n11271), .IN2(n11852), .IN3(n14304), .IN4(n11847), .Q(
        n11251) );
  OA22X1 U4616 ( .IN1(n11271), .IN2(n11851), .IN3(n14304), .IN4(n11846), .Q(
        n11255) );
  XOR2X1 U4619 ( .IN1(n14940), .IN2(n11277), .Q(n11276) );
  AO22X1 U4624 ( .IN1(\fadd_0_0_0_0_10/U24/DATA2_1 ), .IN2(n14963), .IN3(
        \fadd_0_0_0_0_10/U24/DATA1_1 ), .IN4(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_dualsubclose/sub_1_root_add_300/carry[6] ), .Q(\fadd_0_0_0_0_10/U24/Z_1 ) );
  AO22X1 U4625 ( .IN1(\fadd_0_0_0_0_10/U24/DATA2_2 ), .IN2(n14963), .IN3(
        \fadd_0_0_0_0_10/U24/DATA1_2 ), .IN4(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_dualsubclose/sub_1_root_add_300/carry[6] ), .Q(\fadd_0_0_0_0_10/U24/Z_2 ) );
  AO21X1 U4626 ( .IN1(n11282), .IN2(n11283), .IN3(n11240), .Q(n11279) );
  XOR2X1 U4627 ( .IN1(\fadd_0_0_0_0_10/U28/Z_4 ), .IN2(n11280), .Q(n11240) );
  OA22X1 U4628 ( .IN1(n11271), .IN2(n11849), .IN3(n14188), .IN4(n11854), .Q(
        n11280) );
  AO22X1 U4629 ( .IN1(n14304), .IN2(n13585), .IN3(n11271), .IN4(n13726), .Q(
        \fadd_0_0_0_0_10/U28/Z_4 ) );
  OR2X1 U4633 ( .IN1(\fadd_0_0_0_0_10/U5/DATA2_3 ), .IN2(
        \fadd_0_0_0_0_10/U5/DATA2_4 ), .Q(n11272) );
  OR4X1 U4634 ( .IN1(n11273), .IN2(n11271), .IN3(\fadd_0_0_0_0_10/U5/DATA1_1 ), 
        .IN4(\fadd_0_0_0_0_10/U5/DATA1_2 ), .Q(n11282) );
  OR2X1 U4635 ( .IN1(\fadd_0_0_0_0_10/U5/DATA1_3 ), .IN2(
        \fadd_0_0_0_0_10/U5/DATA1_4 ), .Q(n11273) );
  OR4X1 U4636 ( .IN1(\fadd_0_0_0_0_10/U24/Z_3 ), .IN2(
        \fadd_0_0_0_0_10/U24/Z_4 ), .IN3(\fadd_0_0_0_0_10/U24/Z_5 ), .IN4(
        n14964), .Q(n11281) );
  OA22X1 U4640 ( .IN1(n11271), .IN2(n11850), .IN3(n14304), .IN4(n11845), .Q(
        n11262) );
  AO22X1 U4641 ( .IN1(\fadd_0_0_0_0_10/U5/DATA1_0 ), .IN2(n14188), .IN3(
        \fadd_0_0_0_0_10/U5/DATA2_0 ), .IN4(n11271), .Q(
        \fadd_0_0_0_0_10/U27/DATA1_0 ) );
  AND2X1 U4644 ( .IN1(n12808), .IN2(n11284), .Q(n11285) );
  OA22X1 U4646 ( .IN1(\fadd_0_0_0_0_10/sub_707/carry[5] ), .IN2(n12809), .IN3(
        n13469), .IN4(n11286), .Q(n11284) );
  AND2X1 U4647 ( .IN1(n12809), .IN2(\fadd_0_0_0_0_10/sub_707/carry[5] ), .Q(
        n11286) );
  AO22X1 U4649 ( .IN1(\fadd_0_0_0_0_10/U24/DATA2_5 ), .IN2(n14963), .IN3(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_dualsubclose/sub_1_root_add_300/carry[6] ), .IN4(\fadd_0_0_0_0_10/U24/DATA1_5 ), .Q(\fadd_0_0_0_0_10/U24/Z_5 ) );
  AO22X1 U4650 ( .IN1(\fadd_0_0_0_0_10/U24/DATA2_4 ), .IN2(n14963), .IN3(
        \fadd_0_0_0_0_10/U24/DATA1_4 ), .IN4(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_dualsubclose/sub_1_root_add_300/carry[6] ), .Q(\fadd_0_0_0_0_10/U24/Z_4 ) );
  AO22X1 U4651 ( .IN1(\fadd_0_0_0_0_10/U24/DATA2_3 ), .IN2(n14963), .IN3(
        \fadd_0_0_0_0_10/U24/DATA1_3 ), .IN4(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_dualsubclose/sub_1_root_add_300/carry[6] ), .Q(\fadd_0_0_0_0_10/U24/Z_3 ) );
  NOR3X0 U4653 ( .IN1(n14929), .IN2(n11494), .IN3(n10411), .QN(
        \fadd_0_0_0_0_1/zerofromclose ) );
  NAND3X0 U4655 ( .IN1(n13680), .IN2(n13488), .IN3(n11291), .QN(n11288) );
  NAND3X0 U4656 ( .IN1(n11292), .IN2(n11293), .IN3(n12839), .QN(n11287) );
  AO222X1 U4661 ( .IN1(\fadd_0_0_0_0_1/fracresultfar0 [1]), .IN2(n14690), 
        .IN3(\fadd_0_0_0_0_1/fracresultfar0 [2]), .IN4(n11297), .IN5(
        \fadd_0_0_0_0_1/fracresultfar0 [0]), .IN6(
        \fadd_0_0_0_0_1/add_859/B[1] ), .Q(n11292) );
  AO22X1 U4662 ( .IN1(n11301), .IN2(
        \fadd_0_0_0_0_1/rightshiftercomponent/ps_d1 [1]), .IN3(n11302), .IN4(
        \fadd_0_0_0_0_1/rightshiftercomponent/ps_d1 [2]), .Q(
        \fadd_0_0_0_0_1/rightshiftercomponent/n389_o ) );
  AO22X1 U4665 ( .IN1(n13649), .IN2(\fadd_0_0_0_0_1/exponentresultclose_d1 [5]), .IN3(\fadd_0_0_0_0_1/exponentresultfar1 [5]), .IN4(n12839), .Q(
        \fadd_0_0_0_0_1/resultbeforeround [9]) );
  AO22X1 U4666 ( .IN1(n13649), .IN2(\fadd_0_0_0_0_1/exponentresultclose_d1 [4]), .IN3(\fadd_0_0_0_0_1/exponentresultfar1 [4]), .IN4(n12839), .Q(
        \fadd_0_0_0_0_1/resultbeforeround [8]) );
  AO22X1 U4667 ( .IN1(n13649), .IN2(\fadd_0_0_0_0_1/exponentresultclose_d1 [3]), .IN3(\fadd_0_0_0_0_1/exponentresultfar1 [3]), .IN4(n12839), .Q(
        \fadd_0_0_0_0_1/resultbeforeround [7]) );
  AO22X1 U4668 ( .IN1(n13649), .IN2(\fadd_0_0_0_0_1/exponentresultclose_d1 [2]), .IN3(\fadd_0_0_0_0_1/exponentresultfar1 [2]), .IN4(n12839), .Q(
        \fadd_0_0_0_0_1/resultbeforeround [6]) );
  AO22X1 U4669 ( .IN1(n13649), .IN2(\fadd_0_0_0_0_1/exponentresultclose_d1 [1]), .IN3(\fadd_0_0_0_0_1/exponentresultfar1 [1]), .IN4(n12839), .Q(
        \fadd_0_0_0_0_1/resultbeforeround [5]) );
  AO22X1 U4670 ( .IN1(n13649), .IN2(\fadd_0_0_0_0_1/exponentresultclose_d1 [0]), .IN3(\fadd_0_0_0_0_1/exponentresultfar1 [0]), .IN4(n12839), .Q(
        \fadd_0_0_0_0_1/resultbeforeround [4]) );
  AO222X1 U4671 ( .IN1(n11291), .IN2(\fadd_0_0_0_0_1/norm/level1_d1[4] ), 
        .IN3(n11304), .IN4(n13701), .IN5(n12839), .IN6(n11306), .Q(
        \fadd_0_0_0_0_1/resultbeforeround [3]) );
  AO222X1 U4672 ( .IN1(\fadd_0_0_0_0_1/fracresultfar0 [5]), .IN2(n14690), 
        .IN3(n11297), .IN4(\fadd_0_0_0_0_1/fracresultfar0 [6]), .IN5(
        \fadd_0_0_0_0_1/fracresultfar0 [4]), .IN6(
        \fadd_0_0_0_0_1/add_859/B[1] ), .Q(n11306) );
  AO222X1 U4673 ( .IN1(n11291), .IN2(n13701), .IN3(n11304), .IN4(n13565), 
        .IN5(n12839), .IN6(n11308), .Q(\fadd_0_0_0_0_1/resultbeforeround [2])
         );
  AO222X1 U4674 ( .IN1(\fadd_0_0_0_0_1/fracresultfar0 [4]), .IN2(n14690), 
        .IN3(\fadd_0_0_0_0_1/fracresultfar0 [5]), .IN4(n11297), .IN5(
        \fadd_0_0_0_0_1/add_859/B[1] ), .IN6(
        \fadd_0_0_0_0_1/fracresultfar0 [3]), .Q(n11308) );
  AO222X1 U4676 ( .IN1(n11291), .IN2(n13565), .IN3(n11304), .IN4(n13488), 
        .IN5(n12839), .IN6(n11309), .Q(\fadd_0_0_0_0_1/resultbeforeround [1])
         );
  AO222X1 U4677 ( .IN1(\fadd_0_0_0_0_1/fracresultfar0 [3]), .IN2(n14690), 
        .IN3(\fadd_0_0_0_0_1/fracresultfar0 [4]), .IN4(n11297), .IN5(
        \fadd_0_0_0_0_1/add_859/B[1] ), .IN6(
        \fadd_0_0_0_0_1/fracresultfar0 [2]), .Q(n11309) );
  AO22X1 U4679 ( .IN1(n13649), .IN2(\fadd_0_0_0_0_1/exponentresultclose_d1 [6]), .IN3(\fadd_0_0_0_0_1/exponentresultfar1 [6]), .IN4(n12839), .Q(
        \fadd_0_0_0_0_1/resultbeforeround [10]) );
  AO222X1 U4680 ( .IN1(n11291), .IN2(n13488), .IN3(n11304), .IN4(n13680), 
        .IN5(n12839), .IN6(n11299), .Q(\fadd_0_0_0_0_1/resultbeforeround [0])
         );
  AO222X1 U4681 ( .IN1(\fadd_0_0_0_0_1/fracresultfar0 [2]), .IN2(n14690), 
        .IN3(\fadd_0_0_0_0_1/fracresultfar0 [3]), .IN4(n11297), .IN5(
        \fadd_0_0_0_0_1/fracresultfar0 [1]), .IN6(
        \fadd_0_0_0_0_1/add_859/B[1] ), .Q(n11299) );
  AND2X1 U4688 ( .IN1(n12851), .IN2(n13649), .Q(n11291) );
  OA221X1 U4690 ( .IN1(n11310), .IN2(n11311), .IN3(n11312), .IN4(n11313), 
        .IN5(n11314), .Q(\fadd_0_0_0_0_1/ressign ) );
  OR4X1 U4695 ( .IN1(\fadd_0_0_0_0_1/fracrcloseymx [2]), .IN2(
        \fadd_0_0_0_0_1/fracrcloseymx [3]), .IN3(
        \fadd_0_0_0_0_1/fracrcloseymx [4]), .IN4(
        \fadd_0_0_0_0_1/fracrcloseymx [5]), .Q(n11312) );
  OR4X1 U4696 ( .IN1(n11317), .IN2(\fadd_0_0_0_0_1/fracrcloseymx [0]), .IN3(
        \fadd_0_0_0_0_1/fracrclosexmy [1]), .IN4(
        \fadd_0_0_0_0_1/fracrclosexmy [2]), .Q(n11311) );
  AO21X1 U4697 ( .IN1(n11318), .IN2(n11319), .IN3(n14678), .Q(n11317) );
  NAND4X0 U4698 ( .IN1(n11321), .IN2(n11322), .IN3(n14686), .IN4(n14685), .QN(
        n11319) );
  NAND4X0 U4699 ( .IN1(n11325), .IN2(n14303), .IN3(n14688), .IN4(n14687), .QN(
        n11318) );
  AO21X1 U4701 ( .IN1(\fadd_0_0_0_0_1/sub_784/B[1] ), .IN2(n14049), .IN3(
        n11330), .Q(\fadd_0_0_0_0_1/norm/level1 [4]) );
  OAI22X1 U4703 ( .IN1(n14929), .IN2(n11485), .IN3(n11331), .IN4(n11885), .QN(
        \fadd_0_0_0_0_1/norm/level1 [3]) );
  OAI22X1 U4704 ( .IN1(n14929), .IN2(n11484), .IN3(n11331), .IN4(n11886), .QN(
        \fadd_0_0_0_0_1/norm/level1 [2]) );
  NOR3X0 U4709 ( .IN1(n13547), .IN2(n8636), .IN3(n11330), .QN(
        \fadd_0_0_0_0_1/sub_784/B[1] ) );
  OAI21X1 U4710 ( .IN1(n10411), .IN2(n11484), .IN3(n11884), .QN(n11330) );
  NAND4X0 U4713 ( .IN1(n11883), .IN2(n11884), .IN3(n11885), .IN4(n11886), .QN(
        n10411) );
  AO22X1 U4714 ( .IN1(n14303), .IN2(n13509), .IN3(n11322), .IN4(n13622), .Q(
        \fadd_0_0_0_0_1/newy_11 ) );
  AO22X1 U4715 ( .IN1(n14303), .IN2(n13502), .IN3(n11322), .IN4(n13889), .Q(
        \fadd_0_0_0_0_1/newy_10 ) );
  AO22X1 U4716 ( .IN1(n14303), .IN2(n5914), .IN3(n11322), .IN4(n5926), .Q(
        \fadd_0_0_0_0_1/newx [8]) );
  AO22X1 U4719 ( .IN1(n14303), .IN2(n5913), .IN3(n11322), .IN4(n5925), .Q(
        \fadd_0_0_0_0_1/newx [7]) );
  AO22X1 U4722 ( .IN1(n14303), .IN2(n5912), .IN3(n11322), .IN4(n5924), .Q(
        \fadd_0_0_0_0_1/newx [6]) );
  AO22X1 U4725 ( .IN1(n14303), .IN2(n5911), .IN3(n11322), .IN4(n5923), .Q(
        \fadd_0_0_0_0_1/newx [5]) );
  AO22X1 U4728 ( .IN1(n14303), .IN2(n5910), .IN3(n11322), .IN4(n5922), .Q(
        \fadd_0_0_0_0_1/newx [4]) );
  AO22X1 U4731 ( .IN1(n14303), .IN2(n13708), .IN3(n11322), .IN4(n13570), .Q(
        \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ) );
  AO22X1 U4734 ( .IN1(n14303), .IN2(n13686), .IN3(n11322), .IN4(n13553), .Q(
        \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ) );
  AO22X1 U4737 ( .IN1(n14303), .IN2(n13665), .IN3(n11322), .IN4(n13528), .Q(
        \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ) );
  AO22X1 U4741 ( .IN1(n14303), .IN2(n13889), .IN3(n11322), .IN4(n13502), .Q(
        \fadd_0_0_0_0_1/newx [10]) );
  AO22X1 U4743 ( .IN1(n14303), .IN2(n13637), .IN3(n11322), .IN4(n13517), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ) );
  XOR2X1 U4746 ( .IN1(n11332), .IN2(n14678), .Q(
        \fadd_0_0_0_0_1/fracyfarxorop [6]) );
  XOR2X1 U4748 ( .IN1(n11335), .IN2(n12702), .Q(
        \fadd_0_0_0_0_1/fracyfarxorop [5]) );
  OA21X1 U4749 ( .IN1(n12699), .IN2(n14680), .IN3(n14675), .Q(n11335) );
  XOR2X1 U4751 ( .IN1(n11338), .IN2(n12702), .Q(
        \fadd_0_0_0_0_1/fracyfarxorop [4]) );
  OA22X1 U4752 ( .IN1(n14677), .IN2(n11339), .IN3(n12699), .IN4(n11340), .Q(
        n11338) );
  AO22X1 U4754 ( .IN1(n11342), .IN2(n14677), .IN3(n11343), .IN4(n12699), .Q(
        \fadd_0_0_0_0_1/fracyfarxorop [3]) );
  XOR2X1 U4755 ( .IN1(n11340), .IN2(n12702), .Q(n11343) );
  AO21X1 U4756 ( .IN1(n14681), .IN2(n11345), .IN3(n14674), .Q(n11340) );
  AO22X1 U4757 ( .IN1(n11347), .IN2(n14677), .IN3(n11342), .IN4(n12699), .Q(
        \fadd_0_0_0_0_1/fracyfarxorop [2]) );
  XOR2X1 U4758 ( .IN1(n14678), .IN2(n11348), .Q(n11342) );
  OA22X1 U4759 ( .IN1(n11341), .IN2(n11349), .IN3(n11350), .IN4(n11337), .Q(
        n11348) );
  AO22X1 U4761 ( .IN1(n11352), .IN2(n14677), .IN3(n11347), .IN4(n12699), .Q(
        \fadd_0_0_0_0_1/fracyfarxorop [1]) );
  XOR2X1 U4762 ( .IN1(n14678), .IN2(n11353), .Q(n11347) );
  OA22X1 U4763 ( .IN1(n11354), .IN2(n11349), .IN3(n14676), .IN4(n11355), .Q(
        n11353) );
  AO22X1 U4765 ( .IN1(n11352), .IN2(n12699), .IN3(n11356), .IN4(n14677), .Q(
        \fadd_0_0_0_0_1/fracyfarxorop [0]) );
  XOR2X1 U4767 ( .IN1(n12700), .IN2(n12702), .Q(n11356) );
  OA22X1 U4768 ( .IN1(n14676), .IN2(n12701), .IN3(n14683), .IN4(n14673), .Q(
        n12700) );
  XOR2X1 U4772 ( .IN1(n14678), .IN2(n11358), .Q(n11352) );
  AOI22X1 U4773 ( .IN1(n14682), .IN2(n14674), .IN3(n11351), .IN4(
        \fadd_0_0_0_0_1/rightshiftercomponent/level2[1] ), .QN(n11358) );
  OA221X1 U4777 ( .IN1(n14685), .IN2(n14303), .IN3(n14687), .IN4(n11322), 
        .IN5(n11357), .Q(n11345) );
  OA221X1 U4781 ( .IN1(n14686), .IN2(n14303), .IN3(n14688), .IN4(n11322), 
        .IN5(n11357), .Q(n11351) );
  OA22X1 U4782 ( .IN1(n14303), .IN2(n11321), .IN3(n11325), .IN4(n11322), .Q(
        n11357) );
  XOR2X1 U4788 ( .IN1(n14679), .IN2(\fadd_0_0_0_0_1/newy_9 ), .Q(n12702) );
  AO22X1 U4789 ( .IN1(n14303), .IN2(n13579), .IN3(n11322), .IN4(n13717), .Q(
        \fadd_0_0_0_0_1/newy_9 ) );
  OA22X1 U4793 ( .IN1(n11322), .IN2(n11665), .IN3(n14303), .IN4(n11676), .Q(
        n11316) );
  AO22X1 U4795 ( .IN1(n14684), .IN2(n14681), .IN3(n14680), .IN4(n11359), .Q(
        \fadd_0_0_0_0_1/fracyclose1 [3]) );
  OA22X1 U4797 ( .IN1(n11322), .IN2(n11670), .IN3(n14303), .IN4(n11659), .Q(
        n11341) );
  AO22X1 U4798 ( .IN1(n14684), .IN2(n14682), .IN3(n14681), .IN4(n11359), .Q(
        \fadd_0_0_0_0_1/fracyclose1 [2]) );
  OA22X1 U4800 ( .IN1(n11322), .IN2(n11669), .IN3(n14303), .IN4(n11658), .Q(
        n11354) );
  AO22X1 U4801 ( .IN1(n14682), .IN2(n11359), .IN3(n14684), .IN4(n14683), .Q(
        \fadd_0_0_0_0_1/fracyclose1 [1]) );
  OA22X1 U4804 ( .IN1(n11322), .IN2(n11668), .IN3(n14303), .IN4(n11657), .Q(
        n11350) );
  OA22X1 U4806 ( .IN1(n11322), .IN2(n11667), .IN3(n14303), .IN4(n11656), .Q(
        n11360) );
  AO22X1 U4808 ( .IN1(\fadd_0_0_0_0_1/exponentdifferenceyx [0]), .IN2(n14303), 
        .IN3(\fadd_0_0_0_0_1/exponentdifferencexy [0]), .IN4(n11322), .Q(
        n11359) );
  OA22X1 U4811 ( .IN1(n11666), .IN2(n11363), .IN3(
        \fadd_0_0_0_0_1/sub_707/carry [5]), .IN4(n13502), .Q(n11362) );
  AO22X1 U4818 ( .IN1(\fadd_0_0_0_0_1/fracrcloseymx [5]), .IN2(n14113), .IN3(
        \fadd_0_0_0_0_1/fracrclosexmy [5]), .IN4(n14641), .Q(
        \fadd_0_0_0_0_1/fracrclose1 [5]) );
  AO22X1 U4819 ( .IN1(\fadd_0_0_0_0_1/fracrcloseymx [4]), .IN2(n14113), .IN3(
        \fadd_0_0_0_0_1/fracrclosexmy [4]), .IN4(n14641), .Q(
        \fadd_0_0_0_0_1/fracrclose1 [4]) );
  AO22X1 U4820 ( .IN1(\fadd_0_0_0_0_1/fracrcloseymx [3]), .IN2(n14113), .IN3(
        \fadd_0_0_0_0_1/fracrclosexmy [3]), .IN4(n14641), .Q(
        \fadd_0_0_0_0_1/fracrclose1 [3]) );
  AO22X1 U4821 ( .IN1(\fadd_0_0_0_0_1/fracrcloseymx [2]), .IN2(n14113), .IN3(
        \fadd_0_0_0_0_1/fracrclosexmy [2]), .IN4(n14641), .Q(
        \fadd_0_0_0_0_1/fracrclose1 [2]) );
  AO22X1 U4822 ( .IN1(\fadd_0_0_0_0_1/fracrcloseymx [1]), .IN2(n14113), .IN3(
        \fadd_0_0_0_0_1/fracrclosexmy [1]), .IN4(n14641), .Q(
        \fadd_0_0_0_0_1/fracrclose1 [1]) );
  AO22X1 U4823 ( .IN1(\fadd_0_0_0_0_1/fracrcloseymx [0]), .IN2(n14113), .IN3(
        \fadd_0_0_0_0_1/fracrcloseymx [0]), .IN4(n14641), .Q(
        \fadd_0_0_0_0_1/fracrclose1 [0]) );
  NOR3X0 U4827 ( .IN1(n14942), .IN2(n11483), .IN3(n11298), .QN(
        \fadd_0_0_0_0_1/cinaddfar ) );
  AND2X1 U4828 ( .IN1(\fadd_0_0_0_0_1/rightshiftercomponent/level1_d2[0] ), 
        .IN2(\fadd_0_0_0_0_1/rightshiftercomponent/ps_d2[0] ), .Q(n11298) );
  NOR3X0 U4830 ( .IN1(n14928), .IN2(n11481), .IN3(n10410), .QN(
        \fadd_0_0_0_0_0/zerofromclose ) );
  NAND3X0 U4832 ( .IN1(n13679), .IN2(n13487), .IN3(n11372), .QN(n11369) );
  NAND3X0 U4833 ( .IN1(n11373), .IN2(n11374), .IN3(n12838), .QN(n11368) );
  AO222X1 U4838 ( .IN1(\fadd_0_0_0_0_0/fracresultfar0 [1]), .IN2(n14669), 
        .IN3(\fadd_0_0_0_0_0/fracresultfar0 [2]), .IN4(n11378), .IN5(
        \fadd_0_0_0_0_0/fracresultfar0 [0]), .IN6(n14224), .Q(n11373) );
  AO22X1 U4839 ( .IN1(n11382), .IN2(
        \fadd_0_0_0_0_0/rightshiftercomponent/ps_d1 [1]), .IN3(n11383), .IN4(
        \fadd_0_0_0_0_0/rightshiftercomponent/ps_d1 [2]), .Q(
        \fadd_0_0_0_0_0/rightshiftercomponent/n389_o ) );
  AO22X1 U4842 ( .IN1(n13648), .IN2(\fadd_0_0_0_0_0/exponentresultclose_d1 [5]), .IN3(\fadd_0_0_0_0_0/exponentresultfar1 [5]), .IN4(n12838), .Q(
        \fadd_0_0_0_0_0/resultbeforeround [9]) );
  AO22X1 U4843 ( .IN1(n13648), .IN2(\fadd_0_0_0_0_0/exponentresultclose_d1 [4]), .IN3(\fadd_0_0_0_0_0/exponentresultfar1 [4]), .IN4(n12838), .Q(
        \fadd_0_0_0_0_0/resultbeforeround [8]) );
  AO22X1 U4844 ( .IN1(n13648), .IN2(\fadd_0_0_0_0_0/exponentresultclose_d1 [3]), .IN3(\fadd_0_0_0_0_0/exponentresultfar1 [3]), .IN4(n12838), .Q(
        \fadd_0_0_0_0_0/resultbeforeround [7]) );
  AO22X1 U4845 ( .IN1(n13648), .IN2(\fadd_0_0_0_0_0/exponentresultclose_d1 [2]), .IN3(\fadd_0_0_0_0_0/exponentresultfar1 [2]), .IN4(n12838), .Q(
        \fadd_0_0_0_0_0/resultbeforeround [6]) );
  AO22X1 U4846 ( .IN1(n13648), .IN2(\fadd_0_0_0_0_0/exponentresultclose_d1 [1]), .IN3(\fadd_0_0_0_0_0/exponentresultfar1 [1]), .IN4(n12838), .Q(
        \fadd_0_0_0_0_0/resultbeforeround [5]) );
  AO22X1 U4847 ( .IN1(n13648), .IN2(\fadd_0_0_0_0_0/exponentresultclose_d1 [0]), .IN3(\fadd_0_0_0_0_0/exponentresultfar1 [0]), .IN4(n12838), .Q(
        \fadd_0_0_0_0_0/resultbeforeround [4]) );
  AO222X1 U4848 ( .IN1(n11372), .IN2(\fadd_0_0_0_0_0/norm/level1_d1[4] ), 
        .IN3(n11385), .IN4(n13700), .IN5(n12838), .IN6(n11387), .Q(
        \fadd_0_0_0_0_0/resultbeforeround [3]) );
  AO222X1 U4849 ( .IN1(\fadd_0_0_0_0_0/fracresultfar0 [5]), .IN2(n14669), 
        .IN3(n11378), .IN4(\fadd_0_0_0_0_0/fracresultfar0 [6]), .IN5(
        \fadd_0_0_0_0_0/fracresultfar0 [4]), .IN6(n14224), .Q(n11387) );
  AO222X1 U4850 ( .IN1(n11372), .IN2(n13700), .IN3(n11385), .IN4(n13564), 
        .IN5(n12838), .IN6(n11389), .Q(\fadd_0_0_0_0_0/resultbeforeround [2])
         );
  AO222X1 U4851 ( .IN1(\fadd_0_0_0_0_0/fracresultfar0 [4]), .IN2(n14669), 
        .IN3(\fadd_0_0_0_0_0/fracresultfar0 [5]), .IN4(n11378), .IN5(n14224), 
        .IN6(\fadd_0_0_0_0_0/fracresultfar0 [3]), .Q(n11389) );
  AO222X1 U4853 ( .IN1(n11372), .IN2(n13564), .IN3(n11385), .IN4(n13487), 
        .IN5(n12838), .IN6(n11390), .Q(\fadd_0_0_0_0_0/resultbeforeround [1])
         );
  AO222X1 U4854 ( .IN1(\fadd_0_0_0_0_0/fracresultfar0 [3]), .IN2(n14669), 
        .IN3(\fadd_0_0_0_0_0/fracresultfar0 [4]), .IN4(n11378), .IN5(n14224), 
        .IN6(\fadd_0_0_0_0_0/fracresultfar0 [2]), .Q(n11390) );
  AO22X1 U4856 ( .IN1(n13648), .IN2(\fadd_0_0_0_0_0/exponentresultclose_d1 [6]), .IN3(\fadd_0_0_0_0_0/exponentresultfar1 [6]), .IN4(n12838), .Q(
        \fadd_0_0_0_0_0/resultbeforeround [10]) );
  AO222X1 U4857 ( .IN1(n11372), .IN2(n13487), .IN3(n11385), .IN4(n13679), 
        .IN5(n12838), .IN6(n11380), .Q(\fadd_0_0_0_0_0/resultbeforeround [0])
         );
  AO222X1 U4858 ( .IN1(\fadd_0_0_0_0_0/fracresultfar0 [2]), .IN2(n14669), 
        .IN3(\fadd_0_0_0_0_0/fracresultfar0 [3]), .IN4(n11378), .IN5(
        \fadd_0_0_0_0_0/fracresultfar0 [1]), .IN6(n14224), .Q(n11380) );
  AND2X1 U4865 ( .IN1(n12849), .IN2(n13648), .Q(n11372) );
  OA221X1 U4867 ( .IN1(n11391), .IN2(n11392), .IN3(n11393), .IN4(n11394), 
        .IN5(n11395), .Q(\fadd_0_0_0_0_0/ressign ) );
  OR4X1 U4872 ( .IN1(\fadd_0_0_0_0_0/fracrcloseymx [2]), .IN2(
        \fadd_0_0_0_0_0/fracrcloseymx [3]), .IN3(
        \fadd_0_0_0_0_0/fracrcloseymx [4]), .IN4(
        \fadd_0_0_0_0_0/fracrcloseymx [5]), .Q(n11393) );
  OR4X1 U4873 ( .IN1(n11398), .IN2(\fadd_0_0_0_0_0/fracrcloseymx [0]), .IN3(
        \fadd_0_0_0_0_0/fracrclosexmy [1]), .IN4(
        \fadd_0_0_0_0_0/fracrclosexmy [2]), .Q(n11392) );
  AO21X1 U4874 ( .IN1(n11399), .IN2(n11400), .IN3(n14657), .Q(n11398) );
  NAND4X0 U4875 ( .IN1(n11402), .IN2(n11403), .IN3(n14665), .IN4(n14664), .QN(
        n11400) );
  NAND4X0 U4876 ( .IN1(n11406), .IN2(n14302), .IN3(n14667), .IN4(n14666), .QN(
        n11399) );
  AO21X1 U4878 ( .IN1(\fadd_0_0_0_0_0/sub_784/B[1] ), .IN2(n14048), .IN3(
        n11411), .Q(\fadd_0_0_0_0_0/norm/level1 [4]) );
  OAI22X1 U4880 ( .IN1(n14928), .IN2(n11472), .IN3(n11412), .IN4(n11881), .QN(
        \fadd_0_0_0_0_0/norm/level1 [3]) );
  OAI22X1 U4881 ( .IN1(n14928), .IN2(n11471), .IN3(n11412), .IN4(n11882), .QN(
        \fadd_0_0_0_0_0/norm/level1 [2]) );
  NOR3X0 U4886 ( .IN1(n13548), .IN2(n8632), .IN3(n11411), .QN(
        \fadd_0_0_0_0_0/sub_784/B[1] ) );
  OAI21X1 U4887 ( .IN1(n10410), .IN2(n11471), .IN3(n11880), .QN(n11411) );
  NAND4X0 U4890 ( .IN1(n11879), .IN2(n11880), .IN3(n11881), .IN4(n11882), .QN(
        n10410) );
  AO22X1 U4891 ( .IN1(n14302), .IN2(n13515), .IN3(n11403), .IN4(n13627), .Q(
        \fadd_0_0_0_0_0/newy_11 ) );
  AO22X1 U4892 ( .IN1(n14302), .IN2(n13506), .IN3(n11403), .IN4(n13894), .Q(
        \fadd_0_0_0_0_0/newy_10 ) );
  AO22X1 U4893 ( .IN1(n14302), .IN2(n5986), .IN3(n11403), .IN4(n5998), .Q(
        \fadd_0_0_0_0_0/newx [8]) );
  AO22X1 U4896 ( .IN1(n14302), .IN2(n5985), .IN3(n11403), .IN4(n5997), .Q(
        \fadd_0_0_0_0_0/newx [7]) );
  AO22X1 U4899 ( .IN1(n14302), .IN2(n5984), .IN3(n11403), .IN4(n5996), .Q(
        \fadd_0_0_0_0_0/newx [6]) );
  AO22X1 U4902 ( .IN1(n14302), .IN2(n5983), .IN3(n11403), .IN4(n5995), .Q(
        \fadd_0_0_0_0_0/newx [5]) );
  AO22X1 U4905 ( .IN1(n14302), .IN2(n5982), .IN3(n11403), .IN4(n5994), .Q(
        \fadd_0_0_0_0_0/newx [4]) );
  AO22X1 U4908 ( .IN1(n14302), .IN2(n13713), .IN3(n11403), .IN4(n13576), .Q(
        \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ) );
  AO22X1 U4911 ( .IN1(n14302), .IN2(n13691), .IN3(n11403), .IN4(n13559), .Q(
        \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ) );
  AO22X1 U4914 ( .IN1(n14302), .IN2(n13670), .IN3(n11403), .IN4(n13534), .Q(
        \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ) );
  AO22X1 U4918 ( .IN1(n14302), .IN2(n13894), .IN3(n11403), .IN4(n13506), .Q(
        \fadd_0_0_0_0_0/newx [10]) );
  AO22X1 U4920 ( .IN1(n14302), .IN2(n13642), .IN3(n11403), .IN4(n13523), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ) );
  XOR2X1 U4923 ( .IN1(n11415), .IN2(n14657), .Q(
        \fadd_0_0_0_0_0/fracyfarxorop [6]) );
  XOR2X1 U4925 ( .IN1(n11418), .IN2(n12694), .Q(
        \fadd_0_0_0_0_0/fracyfarxorop [5]) );
  OA21X1 U4926 ( .IN1(n12691), .IN2(n14659), .IN3(n14654), .Q(n11418) );
  XOR2X1 U4928 ( .IN1(n11421), .IN2(n12694), .Q(
        \fadd_0_0_0_0_0/fracyfarxorop [4]) );
  OA22X1 U4929 ( .IN1(n14656), .IN2(n11422), .IN3(n12691), .IN4(n11423), .Q(
        n11421) );
  AO22X1 U4931 ( .IN1(n11425), .IN2(n14656), .IN3(n11426), .IN4(n12691), .Q(
        \fadd_0_0_0_0_0/fracyfarxorop [3]) );
  XOR2X1 U4932 ( .IN1(n11423), .IN2(n12694), .Q(n11426) );
  AO21X1 U4933 ( .IN1(n14660), .IN2(n11428), .IN3(n14653), .Q(n11423) );
  AO22X1 U4934 ( .IN1(n11430), .IN2(n14656), .IN3(n11425), .IN4(n12691), .Q(
        \fadd_0_0_0_0_0/fracyfarxorop [2]) );
  XOR2X1 U4935 ( .IN1(n14657), .IN2(n11431), .Q(n11425) );
  OA22X1 U4936 ( .IN1(n11424), .IN2(n11432), .IN3(n11433), .IN4(n11420), .Q(
        n11431) );
  AO22X1 U4938 ( .IN1(n11435), .IN2(n14656), .IN3(n11430), .IN4(n12691), .Q(
        \fadd_0_0_0_0_0/fracyfarxorop [1]) );
  XOR2X1 U4939 ( .IN1(n14657), .IN2(n11436), .Q(n11430) );
  OA22X1 U4940 ( .IN1(n11437), .IN2(n11432), .IN3(n14655), .IN4(n11438), .Q(
        n11436) );
  AO22X1 U4942 ( .IN1(n11435), .IN2(n12691), .IN3(n11439), .IN4(n14656), .Q(
        \fadd_0_0_0_0_0/fracyfarxorop [0]) );
  XOR2X1 U4944 ( .IN1(n12692), .IN2(n12694), .Q(n11439) );
  OA22X1 U4945 ( .IN1(n14655), .IN2(n12693), .IN3(n14662), .IN4(n14652), .Q(
        n12692) );
  XOR2X1 U4949 ( .IN1(n14657), .IN2(n11441), .Q(n11435) );
  AOI22X1 U4950 ( .IN1(n14661), .IN2(n14653), .IN3(n11434), .IN4(
        \fadd_0_0_0_0_0/rightshiftercomponent/level2[1] ), .QN(n11441) );
  OA221X1 U4954 ( .IN1(n14664), .IN2(n14302), .IN3(n14666), .IN4(n11403), 
        .IN5(n11440), .Q(n11428) );
  OA221X1 U4958 ( .IN1(n14665), .IN2(n14302), .IN3(n14667), .IN4(n11403), 
        .IN5(n11440), .Q(n11434) );
  OA22X1 U4959 ( .IN1(n14302), .IN2(n11402), .IN3(n11406), .IN4(n11403), .Q(
        n11440) );
  XOR2X1 U4965 ( .IN1(n14658), .IN2(\fadd_0_0_0_0_0/newy_9 ), .Q(n12694) );
  OAI22X1 U4966 ( .IN1(n11403), .IN2(n11823), .IN3(n14302), .IN4(n11812), .QN(
        \fadd_0_0_0_0_0/newy_9 ) );
  OA22X1 U4968 ( .IN1(n11403), .IN2(n11812), .IN3(n14302), .IN4(n11823), .Q(
        n11397) );
  AO22X1 U4970 ( .IN1(n14663), .IN2(n14660), .IN3(n14659), .IN4(n11442), .Q(
        \fadd_0_0_0_0_0/fracyclose1 [3]) );
  OA22X1 U4972 ( .IN1(n11403), .IN2(n11817), .IN3(n14302), .IN4(n11806), .Q(
        n11424) );
  AO22X1 U4973 ( .IN1(n14663), .IN2(n14661), .IN3(n14660), .IN4(n11442), .Q(
        \fadd_0_0_0_0_0/fracyclose1 [2]) );
  OA22X1 U4975 ( .IN1(n11403), .IN2(n11816), .IN3(n14302), .IN4(n11805), .Q(
        n11437) );
  AO22X1 U4976 ( .IN1(n14661), .IN2(n11442), .IN3(n14663), .IN4(n14662), .Q(
        \fadd_0_0_0_0_0/fracyclose1 [1]) );
  OA22X1 U4979 ( .IN1(n11403), .IN2(n11815), .IN3(n14302), .IN4(n11804), .Q(
        n11433) );
  OA22X1 U4981 ( .IN1(n11403), .IN2(n11814), .IN3(n14302), .IN4(n11803), .Q(
        n11443) );
  AO22X1 U4983 ( .IN1(\fadd_0_0_0_0_0/exponentdifferenceyx [0]), .IN2(n14302), 
        .IN3(\fadd_0_0_0_0_0/exponentdifferencexy [0]), .IN4(n11403), .Q(
        n11442) );
  OA22X1 U4986 ( .IN1(n11813), .IN2(n11446), .IN3(
        \fadd_0_0_0_0_0/sub_707/carry [5]), .IN4(n13506), .Q(n11445) );
  AO22X1 U4993 ( .IN1(\fadd_0_0_0_0_0/fracrcloseymx [5]), .IN2(n14109), .IN3(
        \fadd_0_0_0_0_0/fracrclosexmy [5]), .IN4(n14648), .Q(
        \fadd_0_0_0_0_0/fracrclose1 [5]) );
  AO22X1 U4994 ( .IN1(\fadd_0_0_0_0_0/fracrcloseymx [4]), .IN2(n14109), .IN3(
        \fadd_0_0_0_0_0/fracrclosexmy [4]), .IN4(n14648), .Q(
        \fadd_0_0_0_0_0/fracrclose1 [4]) );
  AO22X1 U4995 ( .IN1(\fadd_0_0_0_0_0/fracrcloseymx [3]), .IN2(n14109), .IN3(
        \fadd_0_0_0_0_0/fracrclosexmy [3]), .IN4(n14648), .Q(
        \fadd_0_0_0_0_0/fracrclose1 [3]) );
  AO22X1 U4996 ( .IN1(\fadd_0_0_0_0_0/fracrcloseymx [2]), .IN2(n14109), .IN3(
        \fadd_0_0_0_0_0/fracrclosexmy [2]), .IN4(n14648), .Q(
        \fadd_0_0_0_0_0/fracrclose1 [2]) );
  AO22X1 U4997 ( .IN1(\fadd_0_0_0_0_0/fracrcloseymx [1]), .IN2(n14109), .IN3(
        \fadd_0_0_0_0_0/fracrclosexmy [1]), .IN4(n14648), .Q(
        \fadd_0_0_0_0_0/fracrclose1 [1]) );
  AO22X1 U4998 ( .IN1(\fadd_0_0_0_0_0/fracrcloseymx [0]), .IN2(n14109), .IN3(
        \fadd_0_0_0_0_0/fracrcloseymx [0]), .IN4(n14648), .Q(
        \fadd_0_0_0_0_0/fracrclose1 [0]) );
  NOR3X0 U5002 ( .IN1(n14958), .IN2(n11470), .IN3(n11379), .QN(
        \fadd_0_0_0_0_0/cinaddfar ) );
  AND2X1 U5003 ( .IN1(\fadd_0_0_0_0_0/rightshiftercomponent/level1_d2[0] ), 
        .IN2(\fadd_0_0_0_0_0/rightshiftercomponent/ps_d2[0] ), .Q(n11379) );
  AND2X1 U5028 ( .IN1(n14440), .IN2(n11935), .Q(\U4/Z_33 ) );
  AND2X1 U5031 ( .IN1(n14440), .IN2(n11936), .Q(\U4/Z_30 ) );
  linear_DW01_add_21 \add_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/add_54  ( 
        .A({1'b0, 1'b1, 
        \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/x_d2 [5:2], 1'b0, 1'b0}), .B(\fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_fracaddfar/y_d2 ), .CI(
        \fadd_0_0_0_0_9/cinaddfar ), .SUM(\fadd_0_0_0_0_9/fracresultfar0 ) );
  linear_DW01_add_23 \add_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/add_54  ( 
        .A({1'b0, 1'b1, 
        \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/x_d2 [5:2], 1'b0, 1'b0}), .B(\fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_fracaddfar/y_d2 ), .CI(
        \fadd_0_0_0_0_8/cinaddfar ), .SUM(\fadd_0_0_0_0_8/fracresultfar0 ) );
  linear_DW01_add_25 \add_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/add_54  ( 
        .A({1'b0, 1'b1, 
        \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/x_d2 [5:2], 1'b0, 1'b0}), .B(\fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_fracaddfar/y_d2 ), .CI(
        \fadd_0_0_0_0_7/cinaddfar ), .SUM(\fadd_0_0_0_0_7/fracresultfar0 ) );
  linear_DW01_add_27 \add_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/add_54  ( 
        .A({1'b0, 1'b1, 
        \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/x_d2 [5:2], 1'b0, 1'b0}), .B(\fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_fracaddfar/y_d2 ), .CI(
        \fadd_0_0_0_0_6/cinaddfar ), .SUM(\fadd_0_0_0_0_6/fracresultfar0 ) );
  linear_DW01_add_29 \add_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/add_54  ( 
        .A({1'b0, 1'b1, 
        \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/x_d2 [5:2], 1'b0, 1'b0}), .B(\fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_fracaddfar/y_d2 ), .CI(
        \fadd_0_0_0_0_5/cinaddfar ), .SUM(\fadd_0_0_0_0_5/fracresultfar0 ) );
  linear_DW01_add_31 \add_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/add_54  ( 
        .A({1'b0, 1'b1, 
        \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/x_d2 [5:2], 1'b0, 1'b0}), .B(\fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_fracaddfar/y_d2 ), .CI(
        \fadd_0_0_0_0_4/cinaddfar ), .SUM(\fadd_0_0_0_0_4/fracresultfar0 ) );
  linear_DW01_add_33 \add_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/add_54  ( 
        .A({1'b0, 1'b1, 
        \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/x_d2 [5:2], 1'b0, 1'b0}), .B(\fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_fracaddfar/y_d2 ), .CI(
        \fadd_0_0_0_0_3/cinaddfar ), .SUM(\fadd_0_0_0_0_3/fracresultfar0 ) );
  linear_DW01_add_35 \add_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/add_54  ( 
        .A({1'b0, 1'b1, 
        \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/x_d2 [5:2], 1'b0, 1'b0}), .B(\fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_fracaddfar/y_d2 ), .CI(
        \fadd_0_0_0_0_2/cinaddfar ), .SUM(\fadd_0_0_0_0_2/fracresultfar0 ) );
  linear_DW01_add_37 \add_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/add_54  ( 
        .A({1'b0, 1'b1, 
        \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/x_d2 [5:2], 1'b0, 1'b0}), .B(\fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_fracaddfar/y_d2 ), .CI(
        \fadd_0_0_0_0_1/cinaddfar ), .SUM(\fadd_0_0_0_0_1/fracresultfar0 ) );
  linear_DW01_add_39 \add_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/add_54  ( 
        .A({1'b0, 1'b1, 
        \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/x_d2 [5:2], 1'b0, 1'b0}), .B(\fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_fracaddfar/y_d2 ), .CI(
        \fadd_0_0_0_0_0/cinaddfar ), .SUM(\fadd_0_0_0_0_0/fracresultfar0 ) );
  linear_DW_mult_uns_0 \fmul_0_0_0_0_0/significandmultiplication/tile_0_mult/mult_18  ( 
        .a({1'b1, n5957, n5956, n5955, n5954}), .b({1'b1, n5945, n5944, n5943, 
        n5942}), .product({\add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/B[1] , 
        \fmul_0_0_0_0_0/sigprod [8:0]}) );
  linear_DW_mult_uns_1 \fmul_0_0_0_0_1/significandmultiplication/tile_0_mult/mult_18  ( 
        .a({1'b1, n5885, n5884, n5883, n5882}), .b({1'b1, n5873, n5872, n5871, 
        n5870}), .product({\add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/B[1] , 
        \fmul_0_0_0_0_1/sigprod [8:0]}) );
  linear_DW_mult_uns_2 \fmul_0_0_0_0_2/significandmultiplication/tile_0_mult/mult_18  ( 
        .a({1'b1, n5813, n5812, n5811, n5810}), .b({1'b1, n5801, n5800, n5799, 
        n5798}), .product({\add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/B[1] , 
        \fmul_0_0_0_0_2/sigprod [8:0]}) );
  linear_DW_mult_uns_3 \fmul_0_0_0_0_3/significandmultiplication/tile_0_mult/mult_18  ( 
        .a({1'b1, n5741, n5740, n5739, n5738}), .b({1'b1, n5729, n5728, n5727, 
        n5726}), .product({\add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/B[1] , 
        \fmul_0_0_0_0_3/sigprod [8:0]}) );
  linear_DW_mult_uns_4 \fmul_0_0_0_0_4/significandmultiplication/tile_0_mult/mult_18  ( 
        .a({1'b1, n5669, n5668, n5667, n5666}), .b({1'b1, n5657, n5656, n5655, 
        n5654}), .product({\add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/B[1] , 
        \fmul_0_0_0_0_4/sigprod [8:0]}) );
  linear_DW_mult_uns_5 \fmul_0_0_0_0_5/significandmultiplication/tile_0_mult/mult_18  ( 
        .a({1'b1, n5597, n5596, n5595, n5594}), .b({1'b1, n5585, n5584, n5583, 
        n5582}), .product({\add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/B[1] , 
        \fmul_0_0_0_0_5/sigprod [8:0]}) );
  linear_DW_mult_uns_6 \fmul_0_0_0_0_6/significandmultiplication/tile_0_mult/mult_18  ( 
        .a({1'b1, n5525, n5524, n5523, n5522}), .b({1'b1, n5513, n5512, n5511, 
        n5510}), .product({\add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/B[1] , 
        \fmul_0_0_0_0_6/sigprod [8:0]}) );
  linear_DW_mult_uns_7 \fmul_0_0_0_0_7/significandmultiplication/tile_0_mult/mult_18  ( 
        .a({1'b1, n5453, n5452, n5451, n5450}), .b({1'b1, n5441, n5440, n5439, 
        n5438}), .product({\add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/B[1] , 
        \fmul_0_0_0_0_7/sigprod [8:0]}) );
  linear_DW_mult_uns_8 \fmul_0_0_0_0_8/significandmultiplication/tile_0_mult/mult_18  ( 
        .a({1'b1, n5381, n5380, n5379, n5378}), .b({1'b1, n5369, n5368, n5367, 
        n5366}), .product({\add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/B[1] , 
        \fmul_0_0_0_0_8/sigprod [8:0]}) );
  linear_DW_mult_uns_9 \fmul_0_0_0_0_9/significandmultiplication/tile_0_mult/mult_18  ( 
        .a({1'b1, n5309, n5308, n5307, n5306}), .b({1'b1, n5297, n5296, n5295, 
        n5294}), .product({\add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/B[1] , 
        \fmul_0_0_0_0_9/sigprod [8:0]}) );
  FADDX1 \fadd_0_0_0_0_9/add_859/U1_1  ( .A(
        \fadd_0_0_0_0_9/exponentresultfar0_d2 [1]), .B(n14233), .CI(
        \fadd_0_0_0_0_9/add_859/carry [1]), .CO(
        \fadd_0_0_0_0_9/add_859/carry [2]), .S(
        \fadd_0_0_0_0_9/exponentresultfar1 [1]) );
  FADDX1 \fadd_0_0_0_0_9/add_859/U1_2  ( .A(
        \fadd_0_0_0_0_9/exponentresultfar0_d2 [2]), .B(n14233), .CI(
        \fadd_0_0_0_0_9/add_859/carry [2]), .CO(
        \fadd_0_0_0_0_9/add_859/carry [3]), .S(
        \fadd_0_0_0_0_9/exponentresultfar1 [2]) );
  FADDX1 \fadd_0_0_0_0_9/add_859/U1_3  ( .A(
        \fadd_0_0_0_0_9/exponentresultfar0_d2 [3]), .B(n14233), .CI(
        \fadd_0_0_0_0_9/add_859/carry [3]), .CO(
        \fadd_0_0_0_0_9/add_859/carry [4]), .S(
        \fadd_0_0_0_0_9/exponentresultfar1 [3]) );
  FADDX1 \fadd_0_0_0_0_9/add_859/U1_4  ( .A(
        \fadd_0_0_0_0_9/exponentresultfar0_d2 [4]), .B(n14233), .CI(
        \fadd_0_0_0_0_9/add_859/carry [4]), .CO(
        \fadd_0_0_0_0_9/add_859/carry [5]), .S(
        \fadd_0_0_0_0_9/exponentresultfar1 [4]) );
  FADDX1 \fadd_0_0_0_0_9/sub_784/U2_1  ( .A(\fadd_0_0_0_0_9/newx_d1 [5]), .B(
        n14937), .CI(\fadd_0_0_0_0_9/sub_784/carry [1]), .CO(
        \fadd_0_0_0_0_9/sub_784/carry [2]), .S(
        \fadd_0_0_0_0_9/exponentresultclose [1]) );
  FADDX1 \fadd_0_0_0_0_9/sub_784/U2_2  ( .A(\fadd_0_0_0_0_9/newx_d1 [6]), .B(
        n10419), .CI(\fadd_0_0_0_0_9/sub_784/carry [2]), .CO(
        \fadd_0_0_0_0_9/sub_784/carry [3]), .S(
        \fadd_0_0_0_0_9/exponentresultclose [2]) );
  FADDX1 \fadd_0_0_0_0_9/sub_710/U2_1  ( .A(n5335), .B(n14638), .CI(
        \fadd_0_0_0_0_9/sub_710/carry [1]), .CO(
        \fadd_0_0_0_0_9/sub_710/carry [2]), .S(
        \fadd_0_0_0_0_9/exponentdifferenceyx [1]) );
  FADDX1 \fadd_0_0_0_0_9/sub_710/U2_2  ( .A(n5336), .B(n14637), .CI(
        \fadd_0_0_0_0_9/sub_710/carry [2]), .CO(
        \fadd_0_0_0_0_9/sub_710/carry [3]), .S(
        \fadd_0_0_0_0_9/exponentdifferenceyx [2]) );
  FADDX1 \fadd_0_0_0_0_9/sub_710/U2_3  ( .A(n5337), .B(n14636), .CI(
        \fadd_0_0_0_0_9/sub_710/carry [3]), .CO(
        \fadd_0_0_0_0_9/sub_710/carry [4]), .S(
        \fadd_0_0_0_0_9/exponentdifferenceyx [3]) );
  FADDX1 \fadd_0_0_0_0_9/sub_707/U2_1  ( .A(n5347), .B(n14633), .CI(
        \fadd_0_0_0_0_9/sub_707/carry [1]), .CO(
        \fadd_0_0_0_0_9/sub_707/carry [2]), .S(
        \fadd_0_0_0_0_9/exponentdifferencexy [1]) );
  FADDX1 \fadd_0_0_0_0_9/sub_707/U2_2  ( .A(n5348), .B(n14632), .CI(
        \fadd_0_0_0_0_9/sub_707/carry [2]), .CO(
        \fadd_0_0_0_0_9/sub_707/carry [3]), .S(
        \fadd_0_0_0_0_9/exponentdifferencexy [2]) );
  FADDX1 \fadd_0_0_0_0_9/sub_707/U2_3  ( .A(n5349), .B(n14631), .CI(
        \fadd_0_0_0_0_9/sub_707/carry [3]), .CO(
        \fadd_0_0_0_0_9/sub_707/carry [4]), .S(
        \fadd_0_0_0_0_9/exponentdifferencexy [3]) );
  FADDX1 \fadd_0_0_0_0_9/sub_707/U2_4  ( .A(n5350), .B(n14630), .CI(
        \fadd_0_0_0_0_9/sub_707/carry [4]), .CO(
        \fadd_0_0_0_0_9/sub_707/carry [5]), .S(
        \fadd_0_0_0_0_9/exponentdifferencexy [4]) );
  FADDX1 \fadd_0_0_0_0_8/add_859/U1_1  ( .A(
        \fadd_0_0_0_0_8/exponentresultfar0_d2 [1]), .B(n14232), .CI(
        \fadd_0_0_0_0_8/add_859/carry [1]), .CO(
        \fadd_0_0_0_0_8/add_859/carry [2]), .S(
        \fadd_0_0_0_0_8/exponentresultfar1 [1]) );
  FADDX1 \fadd_0_0_0_0_8/add_859/U1_2  ( .A(
        \fadd_0_0_0_0_8/exponentresultfar0_d2 [2]), .B(n14232), .CI(
        \fadd_0_0_0_0_8/add_859/carry [2]), .CO(
        \fadd_0_0_0_0_8/add_859/carry [3]), .S(
        \fadd_0_0_0_0_8/exponentresultfar1 [2]) );
  FADDX1 \fadd_0_0_0_0_8/add_859/U1_3  ( .A(
        \fadd_0_0_0_0_8/exponentresultfar0_d2 [3]), .B(n14232), .CI(
        \fadd_0_0_0_0_8/add_859/carry [3]), .CO(
        \fadd_0_0_0_0_8/add_859/carry [4]), .S(
        \fadd_0_0_0_0_8/exponentresultfar1 [3]) );
  FADDX1 \fadd_0_0_0_0_8/add_859/U1_4  ( .A(
        \fadd_0_0_0_0_8/exponentresultfar0_d2 [4]), .B(n14232), .CI(
        \fadd_0_0_0_0_8/add_859/carry [4]), .CO(
        \fadd_0_0_0_0_8/add_859/carry [5]), .S(
        \fadd_0_0_0_0_8/exponentresultfar1 [4]) );
  FADDX1 \fadd_0_0_0_0_8/sub_784/U2_1  ( .A(\fadd_0_0_0_0_8/newx_d1 [5]), .B(
        n14936), .CI(\fadd_0_0_0_0_8/sub_784/carry [1]), .CO(
        \fadd_0_0_0_0_8/sub_784/carry [2]), .S(
        \fadd_0_0_0_0_8/exponentresultclose [1]) );
  FADDX1 \fadd_0_0_0_0_8/sub_784/U2_2  ( .A(\fadd_0_0_0_0_8/newx_d1 [6]), .B(
        n10418), .CI(\fadd_0_0_0_0_8/sub_784/carry [2]), .CO(
        \fadd_0_0_0_0_8/sub_784/carry [3]), .S(
        \fadd_0_0_0_0_8/exponentresultclose [2]) );
  FADDX1 \fadd_0_0_0_0_8/sub_710/U2_1  ( .A(n5407), .B(n14627), .CI(
        \fadd_0_0_0_0_8/sub_710/carry [1]), .CO(
        \fadd_0_0_0_0_8/sub_710/carry [2]), .S(
        \fadd_0_0_0_0_8/exponentdifferenceyx [1]) );
  FADDX1 \fadd_0_0_0_0_8/sub_710/U2_2  ( .A(n5408), .B(n14626), .CI(
        \fadd_0_0_0_0_8/sub_710/carry [2]), .CO(
        \fadd_0_0_0_0_8/sub_710/carry [3]), .S(
        \fadd_0_0_0_0_8/exponentdifferenceyx [2]) );
  FADDX1 \fadd_0_0_0_0_8/sub_710/U2_3  ( .A(n5409), .B(n14625), .CI(
        \fadd_0_0_0_0_8/sub_710/carry [3]), .CO(
        \fadd_0_0_0_0_8/sub_710/carry [4]), .S(
        \fadd_0_0_0_0_8/exponentdifferenceyx [3]) );
  FADDX1 \fadd_0_0_0_0_8/sub_707/U2_1  ( .A(n5419), .B(n14622), .CI(
        \fadd_0_0_0_0_8/sub_707/carry [1]), .CO(
        \fadd_0_0_0_0_8/sub_707/carry [2]), .S(
        \fadd_0_0_0_0_8/exponentdifferencexy [1]) );
  FADDX1 \fadd_0_0_0_0_8/sub_707/U2_2  ( .A(n5420), .B(n14621), .CI(
        \fadd_0_0_0_0_8/sub_707/carry [2]), .CO(
        \fadd_0_0_0_0_8/sub_707/carry [3]), .S(
        \fadd_0_0_0_0_8/exponentdifferencexy [2]) );
  FADDX1 \fadd_0_0_0_0_8/sub_707/U2_3  ( .A(n5421), .B(n14620), .CI(
        \fadd_0_0_0_0_8/sub_707/carry [3]), .CO(
        \fadd_0_0_0_0_8/sub_707/carry [4]), .S(
        \fadd_0_0_0_0_8/exponentdifferencexy [3]) );
  FADDX1 \fadd_0_0_0_0_8/sub_707/U2_4  ( .A(n5422), .B(n14619), .CI(
        \fadd_0_0_0_0_8/sub_707/carry [4]), .CO(
        \fadd_0_0_0_0_8/sub_707/carry [5]), .S(
        \fadd_0_0_0_0_8/exponentdifferencexy [4]) );
  FADDX1 \fadd_0_0_0_0_7/add_859/U1_1  ( .A(
        \fadd_0_0_0_0_7/exponentresultfar0_d2 [1]), .B(
        \fadd_0_0_0_0_7/add_859/B[1] ), .CI(\fadd_0_0_0_0_7/add_859/carry [1]), 
        .CO(\fadd_0_0_0_0_7/add_859/carry [2]), .S(
        \fadd_0_0_0_0_7/exponentresultfar1 [1]) );
  FADDX1 \fadd_0_0_0_0_7/add_859/U1_2  ( .A(
        \fadd_0_0_0_0_7/exponentresultfar0_d2 [2]), .B(
        \fadd_0_0_0_0_7/add_859/B[1] ), .CI(\fadd_0_0_0_0_7/add_859/carry [2]), 
        .CO(\fadd_0_0_0_0_7/add_859/carry [3]), .S(
        \fadd_0_0_0_0_7/exponentresultfar1 [2]) );
  FADDX1 \fadd_0_0_0_0_7/add_859/U1_3  ( .A(
        \fadd_0_0_0_0_7/exponentresultfar0_d2 [3]), .B(
        \fadd_0_0_0_0_7/add_859/B[1] ), .CI(\fadd_0_0_0_0_7/add_859/carry [3]), 
        .CO(\fadd_0_0_0_0_7/add_859/carry [4]), .S(
        \fadd_0_0_0_0_7/exponentresultfar1 [3]) );
  FADDX1 \fadd_0_0_0_0_7/add_859/U1_4  ( .A(
        \fadd_0_0_0_0_7/exponentresultfar0_d2 [4]), .B(n14231), .CI(
        \fadd_0_0_0_0_7/add_859/carry [4]), .CO(
        \fadd_0_0_0_0_7/add_859/carry [5]), .S(
        \fadd_0_0_0_0_7/exponentresultfar1 [4]) );
  FADDX1 \fadd_0_0_0_0_7/sub_784/U2_1  ( .A(\fadd_0_0_0_0_7/newx_d1 [5]), .B(
        n14935), .CI(\fadd_0_0_0_0_7/sub_784/carry [1]), .CO(
        \fadd_0_0_0_0_7/sub_784/carry [2]), .S(
        \fadd_0_0_0_0_7/exponentresultclose [1]) );
  FADDX1 \fadd_0_0_0_0_7/sub_784/U2_2  ( .A(\fadd_0_0_0_0_7/newx_d1 [6]), .B(
        n10417), .CI(\fadd_0_0_0_0_7/sub_784/carry [2]), .CO(
        \fadd_0_0_0_0_7/sub_784/carry [3]), .S(
        \fadd_0_0_0_0_7/exponentresultclose [2]) );
  FADDX1 \fadd_0_0_0_0_7/sub_710/U2_1  ( .A(n5479), .B(n14616), .CI(
        \fadd_0_0_0_0_7/sub_710/carry [1]), .CO(
        \fadd_0_0_0_0_7/sub_710/carry [2]), .S(
        \fadd_0_0_0_0_7/exponentdifferenceyx [1]) );
  FADDX1 \fadd_0_0_0_0_7/sub_710/U2_2  ( .A(n5480), .B(n14615), .CI(
        \fadd_0_0_0_0_7/sub_710/carry [2]), .CO(
        \fadd_0_0_0_0_7/sub_710/carry [3]), .S(
        \fadd_0_0_0_0_7/exponentdifferenceyx [2]) );
  FADDX1 \fadd_0_0_0_0_7/sub_710/U2_3  ( .A(n5481), .B(n14614), .CI(
        \fadd_0_0_0_0_7/sub_710/carry [3]), .CO(
        \fadd_0_0_0_0_7/sub_710/carry [4]), .S(
        \fadd_0_0_0_0_7/exponentdifferenceyx [3]) );
  FADDX1 \fadd_0_0_0_0_7/sub_707/U2_1  ( .A(n5491), .B(n14611), .CI(
        \fadd_0_0_0_0_7/sub_707/carry [1]), .CO(
        \fadd_0_0_0_0_7/sub_707/carry [2]), .S(
        \fadd_0_0_0_0_7/exponentdifferencexy [1]) );
  FADDX1 \fadd_0_0_0_0_7/sub_707/U2_2  ( .A(n5492), .B(n14610), .CI(
        \fadd_0_0_0_0_7/sub_707/carry [2]), .CO(
        \fadd_0_0_0_0_7/sub_707/carry [3]), .S(
        \fadd_0_0_0_0_7/exponentdifferencexy [2]) );
  FADDX1 \fadd_0_0_0_0_7/sub_707/U2_3  ( .A(n5493), .B(n14609), .CI(
        \fadd_0_0_0_0_7/sub_707/carry [3]), .CO(
        \fadd_0_0_0_0_7/sub_707/carry [4]), .S(
        \fadd_0_0_0_0_7/exponentdifferencexy [3]) );
  FADDX1 \fadd_0_0_0_0_7/sub_707/U2_4  ( .A(n5494), .B(n14608), .CI(
        \fadd_0_0_0_0_7/sub_707/carry [4]), .CO(
        \fadd_0_0_0_0_7/sub_707/carry [5]), .S(
        \fadd_0_0_0_0_7/exponentdifferencexy [4]) );
  FADDX1 \fadd_0_0_0_0_6/add_859/U1_1  ( .A(
        \fadd_0_0_0_0_6/exponentresultfar0_d2 [1]), .B(n14230), .CI(
        \fadd_0_0_0_0_6/add_859/carry [1]), .CO(
        \fadd_0_0_0_0_6/add_859/carry [2]), .S(
        \fadd_0_0_0_0_6/exponentresultfar1 [1]) );
  FADDX1 \fadd_0_0_0_0_6/add_859/U1_2  ( .A(
        \fadd_0_0_0_0_6/exponentresultfar0_d2 [2]), .B(n14230), .CI(
        \fadd_0_0_0_0_6/add_859/carry [2]), .CO(
        \fadd_0_0_0_0_6/add_859/carry [3]), .S(
        \fadd_0_0_0_0_6/exponentresultfar1 [2]) );
  FADDX1 \fadd_0_0_0_0_6/add_859/U1_3  ( .A(
        \fadd_0_0_0_0_6/exponentresultfar0_d2 [3]), .B(n14230), .CI(
        \fadd_0_0_0_0_6/add_859/carry [3]), .CO(
        \fadd_0_0_0_0_6/add_859/carry [4]), .S(
        \fadd_0_0_0_0_6/exponentresultfar1 [3]) );
  FADDX1 \fadd_0_0_0_0_6/add_859/U1_4  ( .A(
        \fadd_0_0_0_0_6/exponentresultfar0_d2 [4]), .B(n14230), .CI(
        \fadd_0_0_0_0_6/add_859/carry [4]), .CO(
        \fadd_0_0_0_0_6/add_859/carry [5]), .S(
        \fadd_0_0_0_0_6/exponentresultfar1 [4]) );
  FADDX1 \fadd_0_0_0_0_6/sub_784/U2_1  ( .A(\fadd_0_0_0_0_6/newx_d1 [5]), .B(
        n14934), .CI(\fadd_0_0_0_0_6/sub_784/carry [1]), .CO(
        \fadd_0_0_0_0_6/sub_784/carry [2]), .S(
        \fadd_0_0_0_0_6/exponentresultclose [1]) );
  FADDX1 \fadd_0_0_0_0_6/sub_784/U2_2  ( .A(\fadd_0_0_0_0_6/newx_d1 [6]), .B(
        n10416), .CI(\fadd_0_0_0_0_6/sub_784/carry [2]), .CO(
        \fadd_0_0_0_0_6/sub_784/carry [3]), .S(
        \fadd_0_0_0_0_6/exponentresultclose [2]) );
  FADDX1 \fadd_0_0_0_0_6/sub_710/U2_1  ( .A(n5551), .B(n14605), .CI(
        \fadd_0_0_0_0_6/sub_710/carry [1]), .CO(
        \fadd_0_0_0_0_6/sub_710/carry [2]), .S(
        \fadd_0_0_0_0_6/exponentdifferenceyx [1]) );
  FADDX1 \fadd_0_0_0_0_6/sub_710/U2_2  ( .A(n5552), .B(n14604), .CI(
        \fadd_0_0_0_0_6/sub_710/carry [2]), .CO(
        \fadd_0_0_0_0_6/sub_710/carry [3]), .S(
        \fadd_0_0_0_0_6/exponentdifferenceyx [2]) );
  FADDX1 \fadd_0_0_0_0_6/sub_710/U2_3  ( .A(n5553), .B(n14603), .CI(
        \fadd_0_0_0_0_6/sub_710/carry [3]), .CO(
        \fadd_0_0_0_0_6/sub_710/carry [4]), .S(
        \fadd_0_0_0_0_6/exponentdifferenceyx [3]) );
  FADDX1 \fadd_0_0_0_0_6/sub_707/U2_1  ( .A(n5563), .B(n14600), .CI(
        \fadd_0_0_0_0_6/sub_707/carry [1]), .CO(
        \fadd_0_0_0_0_6/sub_707/carry [2]), .S(
        \fadd_0_0_0_0_6/exponentdifferencexy [1]) );
  FADDX1 \fadd_0_0_0_0_6/sub_707/U2_2  ( .A(n5564), .B(n14599), .CI(
        \fadd_0_0_0_0_6/sub_707/carry [2]), .CO(
        \fadd_0_0_0_0_6/sub_707/carry [3]), .S(
        \fadd_0_0_0_0_6/exponentdifferencexy [2]) );
  FADDX1 \fadd_0_0_0_0_6/sub_707/U2_3  ( .A(n5565), .B(n14598), .CI(
        \fadd_0_0_0_0_6/sub_707/carry [3]), .CO(
        \fadd_0_0_0_0_6/sub_707/carry [4]), .S(
        \fadd_0_0_0_0_6/exponentdifferencexy [3]) );
  FADDX1 \fadd_0_0_0_0_6/sub_707/U2_4  ( .A(n5566), .B(n14597), .CI(
        \fadd_0_0_0_0_6/sub_707/carry [4]), .CO(
        \fadd_0_0_0_0_6/sub_707/carry [5]), .S(
        \fadd_0_0_0_0_6/exponentdifferencexy [4]) );
  FADDX1 \fadd_0_0_0_0_5/add_859/U1_1  ( .A(
        \fadd_0_0_0_0_5/exponentresultfar0_d2 [1]), .B(
        \fadd_0_0_0_0_5/add_859/B[1] ), .CI(\fadd_0_0_0_0_5/add_859/carry [1]), 
        .CO(\fadd_0_0_0_0_5/add_859/carry [2]), .S(
        \fadd_0_0_0_0_5/exponentresultfar1 [1]) );
  FADDX1 \fadd_0_0_0_0_5/add_859/U1_2  ( .A(
        \fadd_0_0_0_0_5/exponentresultfar0_d2 [2]), .B(
        \fadd_0_0_0_0_5/add_859/B[1] ), .CI(\fadd_0_0_0_0_5/add_859/carry [2]), 
        .CO(\fadd_0_0_0_0_5/add_859/carry [3]), .S(
        \fadd_0_0_0_0_5/exponentresultfar1 [2]) );
  FADDX1 \fadd_0_0_0_0_5/add_859/U1_3  ( .A(
        \fadd_0_0_0_0_5/exponentresultfar0_d2 [3]), .B(
        \fadd_0_0_0_0_5/add_859/B[1] ), .CI(\fadd_0_0_0_0_5/add_859/carry [3]), 
        .CO(\fadd_0_0_0_0_5/add_859/carry [4]), .S(
        \fadd_0_0_0_0_5/exponentresultfar1 [3]) );
  FADDX1 \fadd_0_0_0_0_5/add_859/U1_4  ( .A(
        \fadd_0_0_0_0_5/exponentresultfar0_d2 [4]), .B(n14229), .CI(
        \fadd_0_0_0_0_5/add_859/carry [4]), .CO(
        \fadd_0_0_0_0_5/add_859/carry [5]), .S(
        \fadd_0_0_0_0_5/exponentresultfar1 [4]) );
  FADDX1 \fadd_0_0_0_0_5/sub_784/U2_1  ( .A(\fadd_0_0_0_0_5/newx_d1 [5]), .B(
        n14933), .CI(\fadd_0_0_0_0_5/sub_784/carry [1]), .CO(
        \fadd_0_0_0_0_5/sub_784/carry [2]), .S(
        \fadd_0_0_0_0_5/exponentresultclose [1]) );
  FADDX1 \fadd_0_0_0_0_5/sub_784/U2_2  ( .A(\fadd_0_0_0_0_5/newx_d1 [6]), .B(
        n10415), .CI(\fadd_0_0_0_0_5/sub_784/carry [2]), .CO(
        \fadd_0_0_0_0_5/sub_784/carry [3]), .S(
        \fadd_0_0_0_0_5/exponentresultclose [2]) );
  FADDX1 \fadd_0_0_0_0_5/sub_710/U2_1  ( .A(n5623), .B(n14594), .CI(
        \fadd_0_0_0_0_5/sub_710/carry [1]), .CO(
        \fadd_0_0_0_0_5/sub_710/carry [2]), .S(
        \fadd_0_0_0_0_5/exponentdifferenceyx [1]) );
  FADDX1 \fadd_0_0_0_0_5/sub_710/U2_2  ( .A(n5624), .B(n14593), .CI(
        \fadd_0_0_0_0_5/sub_710/carry [2]), .CO(
        \fadd_0_0_0_0_5/sub_710/carry [3]), .S(
        \fadd_0_0_0_0_5/exponentdifferenceyx [2]) );
  FADDX1 \fadd_0_0_0_0_5/sub_710/U2_3  ( .A(n5625), .B(n14592), .CI(
        \fadd_0_0_0_0_5/sub_710/carry [3]), .CO(
        \fadd_0_0_0_0_5/sub_710/carry [4]), .S(
        \fadd_0_0_0_0_5/exponentdifferenceyx [3]) );
  FADDX1 \fadd_0_0_0_0_5/sub_707/U2_1  ( .A(n5635), .B(n14589), .CI(
        \fadd_0_0_0_0_5/sub_707/carry [1]), .CO(
        \fadd_0_0_0_0_5/sub_707/carry [2]), .S(
        \fadd_0_0_0_0_5/exponentdifferencexy [1]) );
  FADDX1 \fadd_0_0_0_0_5/sub_707/U2_2  ( .A(n5636), .B(n14588), .CI(
        \fadd_0_0_0_0_5/sub_707/carry [2]), .CO(
        \fadd_0_0_0_0_5/sub_707/carry [3]), .S(
        \fadd_0_0_0_0_5/exponentdifferencexy [2]) );
  FADDX1 \fadd_0_0_0_0_5/sub_707/U2_3  ( .A(n5637), .B(n14587), .CI(
        \fadd_0_0_0_0_5/sub_707/carry [3]), .CO(
        \fadd_0_0_0_0_5/sub_707/carry [4]), .S(
        \fadd_0_0_0_0_5/exponentdifferencexy [3]) );
  FADDX1 \fadd_0_0_0_0_5/sub_707/U2_4  ( .A(n5638), .B(n14586), .CI(
        \fadd_0_0_0_0_5/sub_707/carry [4]), .CO(
        \fadd_0_0_0_0_5/sub_707/carry [5]), .S(
        \fadd_0_0_0_0_5/exponentdifferencexy [4]) );
  FADDX1 \fadd_0_0_0_0_4/add_859/U1_1  ( .A(
        \fadd_0_0_0_0_4/exponentresultfar0_d2 [1]), .B(
        \fadd_0_0_0_0_4/add_859/B[1] ), .CI(\fadd_0_0_0_0_4/add_859/carry [1]), 
        .CO(\fadd_0_0_0_0_4/add_859/carry [2]), .S(
        \fadd_0_0_0_0_4/exponentresultfar1 [1]) );
  FADDX1 \fadd_0_0_0_0_4/add_859/U1_2  ( .A(
        \fadd_0_0_0_0_4/exponentresultfar0_d2 [2]), .B(
        \fadd_0_0_0_0_4/add_859/B[1] ), .CI(\fadd_0_0_0_0_4/add_859/carry [2]), 
        .CO(\fadd_0_0_0_0_4/add_859/carry [3]), .S(
        \fadd_0_0_0_0_4/exponentresultfar1 [2]) );
  FADDX1 \fadd_0_0_0_0_4/add_859/U1_3  ( .A(
        \fadd_0_0_0_0_4/exponentresultfar0_d2 [3]), .B(
        \fadd_0_0_0_0_4/add_859/B[1] ), .CI(\fadd_0_0_0_0_4/add_859/carry [3]), 
        .CO(\fadd_0_0_0_0_4/add_859/carry [4]), .S(
        \fadd_0_0_0_0_4/exponentresultfar1 [3]) );
  FADDX1 \fadd_0_0_0_0_4/add_859/U1_4  ( .A(
        \fadd_0_0_0_0_4/exponentresultfar0_d2 [4]), .B(n14228), .CI(
        \fadd_0_0_0_0_4/add_859/carry [4]), .CO(
        \fadd_0_0_0_0_4/add_859/carry [5]), .S(
        \fadd_0_0_0_0_4/exponentresultfar1 [4]) );
  FADDX1 \fadd_0_0_0_0_4/sub_784/U2_1  ( .A(\fadd_0_0_0_0_4/newx_d1 [5]), .B(
        n14932), .CI(\fadd_0_0_0_0_4/sub_784/carry [1]), .CO(
        \fadd_0_0_0_0_4/sub_784/carry [2]), .S(
        \fadd_0_0_0_0_4/exponentresultclose [1]) );
  FADDX1 \fadd_0_0_0_0_4/sub_784/U2_2  ( .A(\fadd_0_0_0_0_4/newx_d1 [6]), .B(
        n10414), .CI(\fadd_0_0_0_0_4/sub_784/carry [2]), .CO(
        \fadd_0_0_0_0_4/sub_784/carry [3]), .S(
        \fadd_0_0_0_0_4/exponentresultclose [2]) );
  FADDX1 \fadd_0_0_0_0_4/sub_710/U2_1  ( .A(n5695), .B(n14583), .CI(
        \fadd_0_0_0_0_4/sub_710/carry [1]), .CO(
        \fadd_0_0_0_0_4/sub_710/carry [2]), .S(
        \fadd_0_0_0_0_4/exponentdifferenceyx [1]) );
  FADDX1 \fadd_0_0_0_0_4/sub_710/U2_2  ( .A(n5696), .B(n14582), .CI(
        \fadd_0_0_0_0_4/sub_710/carry [2]), .CO(
        \fadd_0_0_0_0_4/sub_710/carry [3]), .S(
        \fadd_0_0_0_0_4/exponentdifferenceyx [2]) );
  FADDX1 \fadd_0_0_0_0_4/sub_710/U2_3  ( .A(n5697), .B(n14581), .CI(
        \fadd_0_0_0_0_4/sub_710/carry [3]), .CO(
        \fadd_0_0_0_0_4/sub_710/carry [4]), .S(
        \fadd_0_0_0_0_4/exponentdifferenceyx [3]) );
  FADDX1 \fadd_0_0_0_0_4/sub_707/U2_1  ( .A(n5707), .B(n14578), .CI(
        \fadd_0_0_0_0_4/sub_707/carry [1]), .CO(
        \fadd_0_0_0_0_4/sub_707/carry [2]), .S(
        \fadd_0_0_0_0_4/exponentdifferencexy [1]) );
  FADDX1 \fadd_0_0_0_0_4/sub_707/U2_2  ( .A(n5708), .B(n14577), .CI(
        \fadd_0_0_0_0_4/sub_707/carry [2]), .CO(
        \fadd_0_0_0_0_4/sub_707/carry [3]), .S(
        \fadd_0_0_0_0_4/exponentdifferencexy [2]) );
  FADDX1 \fadd_0_0_0_0_4/sub_707/U2_3  ( .A(n5709), .B(n14576), .CI(
        \fadd_0_0_0_0_4/sub_707/carry [3]), .CO(
        \fadd_0_0_0_0_4/sub_707/carry [4]), .S(
        \fadd_0_0_0_0_4/exponentdifferencexy [3]) );
  FADDX1 \fadd_0_0_0_0_4/sub_707/U2_4  ( .A(n5710), .B(n14575), .CI(
        \fadd_0_0_0_0_4/sub_707/carry [4]), .CO(
        \fadd_0_0_0_0_4/sub_707/carry [5]), .S(
        \fadd_0_0_0_0_4/exponentdifferencexy [4]) );
  FADDX1 \fadd_0_0_0_0_3/add_859/U1_1  ( .A(
        \fadd_0_0_0_0_3/exponentresultfar0_d2 [1]), .B(
        \fadd_0_0_0_0_3/add_859/B[1] ), .CI(\fadd_0_0_0_0_3/add_859/carry [1]), 
        .CO(\fadd_0_0_0_0_3/add_859/carry [2]), .S(
        \fadd_0_0_0_0_3/exponentresultfar1 [1]) );
  FADDX1 \fadd_0_0_0_0_3/add_859/U1_2  ( .A(
        \fadd_0_0_0_0_3/exponentresultfar0_d2 [2]), .B(
        \fadd_0_0_0_0_3/add_859/B[1] ), .CI(\fadd_0_0_0_0_3/add_859/carry [2]), 
        .CO(\fadd_0_0_0_0_3/add_859/carry [3]), .S(
        \fadd_0_0_0_0_3/exponentresultfar1 [2]) );
  FADDX1 \fadd_0_0_0_0_3/add_859/U1_3  ( .A(
        \fadd_0_0_0_0_3/exponentresultfar0_d2 [3]), .B(
        \fadd_0_0_0_0_3/add_859/B[1] ), .CI(\fadd_0_0_0_0_3/add_859/carry [3]), 
        .CO(\fadd_0_0_0_0_3/add_859/carry [4]), .S(
        \fadd_0_0_0_0_3/exponentresultfar1 [3]) );
  FADDX1 \fadd_0_0_0_0_3/add_859/U1_4  ( .A(
        \fadd_0_0_0_0_3/exponentresultfar0_d2 [4]), .B(n14227), .CI(
        \fadd_0_0_0_0_3/add_859/carry [4]), .CO(
        \fadd_0_0_0_0_3/add_859/carry [5]), .S(
        \fadd_0_0_0_0_3/exponentresultfar1 [4]) );
  FADDX1 \fadd_0_0_0_0_3/sub_784/U2_1  ( .A(\fadd_0_0_0_0_3/newx_d1 [5]), .B(
        n14931), .CI(\fadd_0_0_0_0_3/sub_784/carry [1]), .CO(
        \fadd_0_0_0_0_3/sub_784/carry [2]), .S(
        \fadd_0_0_0_0_3/exponentresultclose [1]) );
  FADDX1 \fadd_0_0_0_0_3/sub_784/U2_2  ( .A(\fadd_0_0_0_0_3/newx_d1 [6]), .B(
        n10413), .CI(\fadd_0_0_0_0_3/sub_784/carry [2]), .CO(
        \fadd_0_0_0_0_3/sub_784/carry [3]), .S(
        \fadd_0_0_0_0_3/exponentresultclose [2]) );
  FADDX1 \fadd_0_0_0_0_3/sub_710/U2_1  ( .A(n5767), .B(n14572), .CI(
        \fadd_0_0_0_0_3/sub_710/carry [1]), .CO(
        \fadd_0_0_0_0_3/sub_710/carry [2]), .S(
        \fadd_0_0_0_0_3/exponentdifferenceyx [1]) );
  FADDX1 \fadd_0_0_0_0_3/sub_710/U2_2  ( .A(n5768), .B(n14571), .CI(
        \fadd_0_0_0_0_3/sub_710/carry [2]), .CO(
        \fadd_0_0_0_0_3/sub_710/carry [3]), .S(
        \fadd_0_0_0_0_3/exponentdifferenceyx [2]) );
  FADDX1 \fadd_0_0_0_0_3/sub_710/U2_3  ( .A(n5769), .B(n14570), .CI(
        \fadd_0_0_0_0_3/sub_710/carry [3]), .CO(
        \fadd_0_0_0_0_3/sub_710/carry [4]), .S(
        \fadd_0_0_0_0_3/exponentdifferenceyx [3]) );
  FADDX1 \fadd_0_0_0_0_3/sub_707/U2_1  ( .A(n5779), .B(n14567), .CI(
        \fadd_0_0_0_0_3/sub_707/carry [1]), .CO(
        \fadd_0_0_0_0_3/sub_707/carry [2]), .S(
        \fadd_0_0_0_0_3/exponentdifferencexy [1]) );
  FADDX1 \fadd_0_0_0_0_3/sub_707/U2_2  ( .A(n5780), .B(n14566), .CI(
        \fadd_0_0_0_0_3/sub_707/carry [2]), .CO(
        \fadd_0_0_0_0_3/sub_707/carry [3]), .S(
        \fadd_0_0_0_0_3/exponentdifferencexy [2]) );
  FADDX1 \fadd_0_0_0_0_3/sub_707/U2_3  ( .A(n5781), .B(n14565), .CI(
        \fadd_0_0_0_0_3/sub_707/carry [3]), .CO(
        \fadd_0_0_0_0_3/sub_707/carry [4]), .S(
        \fadd_0_0_0_0_3/exponentdifferencexy [3]) );
  FADDX1 \fadd_0_0_0_0_3/sub_707/U2_4  ( .A(n5782), .B(n14564), .CI(
        \fadd_0_0_0_0_3/sub_707/carry [4]), .CO(
        \fadd_0_0_0_0_3/sub_707/carry [5]), .S(
        \fadd_0_0_0_0_3/exponentdifferencexy [4]) );
  FADDX1 \fadd_0_0_0_0_2/add_859/U1_1  ( .A(
        \fadd_0_0_0_0_2/exponentresultfar0_d2 [1]), .B(
        \fadd_0_0_0_0_2/add_859/B[1] ), .CI(\fadd_0_0_0_0_2/add_859/carry [1]), 
        .CO(\fadd_0_0_0_0_2/add_859/carry [2]), .S(
        \fadd_0_0_0_0_2/exponentresultfar1 [1]) );
  FADDX1 \fadd_0_0_0_0_2/add_859/U1_2  ( .A(
        \fadd_0_0_0_0_2/exponentresultfar0_d2 [2]), .B(
        \fadd_0_0_0_0_2/add_859/B[1] ), .CI(\fadd_0_0_0_0_2/add_859/carry [2]), 
        .CO(\fadd_0_0_0_0_2/add_859/carry [3]), .S(
        \fadd_0_0_0_0_2/exponentresultfar1 [2]) );
  FADDX1 \fadd_0_0_0_0_2/add_859/U1_3  ( .A(
        \fadd_0_0_0_0_2/exponentresultfar0_d2 [3]), .B(
        \fadd_0_0_0_0_2/add_859/B[1] ), .CI(\fadd_0_0_0_0_2/add_859/carry [3]), 
        .CO(\fadd_0_0_0_0_2/add_859/carry [4]), .S(
        \fadd_0_0_0_0_2/exponentresultfar1 [3]) );
  FADDX1 \fadd_0_0_0_0_2/add_859/U1_4  ( .A(
        \fadd_0_0_0_0_2/exponentresultfar0_d2 [4]), .B(n14226), .CI(
        \fadd_0_0_0_0_2/add_859/carry [4]), .CO(
        \fadd_0_0_0_0_2/add_859/carry [5]), .S(
        \fadd_0_0_0_0_2/exponentresultfar1 [4]) );
  FADDX1 \fadd_0_0_0_0_2/sub_784/U2_1  ( .A(\fadd_0_0_0_0_2/newx_d1 [5]), .B(
        n14930), .CI(\fadd_0_0_0_0_2/sub_784/carry [1]), .CO(
        \fadd_0_0_0_0_2/sub_784/carry [2]), .S(
        \fadd_0_0_0_0_2/exponentresultclose [1]) );
  FADDX1 \fadd_0_0_0_0_2/sub_784/U2_2  ( .A(\fadd_0_0_0_0_2/newx_d1 [6]), .B(
        n10412), .CI(\fadd_0_0_0_0_2/sub_784/carry [2]), .CO(
        \fadd_0_0_0_0_2/sub_784/carry [3]), .S(
        \fadd_0_0_0_0_2/exponentresultclose [2]) );
  FADDX1 \fadd_0_0_0_0_2/sub_710/U2_1  ( .A(n5839), .B(n14560), .CI(
        \fadd_0_0_0_0_2/sub_710/carry [1]), .CO(
        \fadd_0_0_0_0_2/sub_710/carry [2]), .S(
        \fadd_0_0_0_0_2/exponentdifferenceyx [1]) );
  FADDX1 \fadd_0_0_0_0_2/sub_710/U2_2  ( .A(n5840), .B(n14559), .CI(
        \fadd_0_0_0_0_2/sub_710/carry [2]), .CO(
        \fadd_0_0_0_0_2/sub_710/carry [3]), .S(
        \fadd_0_0_0_0_2/exponentdifferenceyx [2]) );
  FADDX1 \fadd_0_0_0_0_2/sub_710/U2_3  ( .A(n5841), .B(n14558), .CI(
        \fadd_0_0_0_0_2/sub_710/carry [3]), .CO(
        \fadd_0_0_0_0_2/sub_710/carry [4]), .S(
        \fadd_0_0_0_0_2/exponentdifferenceyx [3]) );
  FADDX1 \fadd_0_0_0_0_2/sub_707/U2_1  ( .A(n5851), .B(n14556), .CI(
        \fadd_0_0_0_0_2/sub_707/carry [1]), .CO(
        \fadd_0_0_0_0_2/sub_707/carry [2]), .S(
        \fadd_0_0_0_0_2/exponentdifferencexy [1]) );
  FADDX1 \fadd_0_0_0_0_2/sub_707/U2_2  ( .A(n5852), .B(n14555), .CI(
        \fadd_0_0_0_0_2/sub_707/carry [2]), .CO(
        \fadd_0_0_0_0_2/sub_707/carry [3]), .S(
        \fadd_0_0_0_0_2/exponentdifferencexy [2]) );
  FADDX1 \fadd_0_0_0_0_2/sub_707/U2_3  ( .A(n5853), .B(n14554), .CI(
        \fadd_0_0_0_0_2/sub_707/carry [3]), .CO(
        \fadd_0_0_0_0_2/sub_707/carry [4]), .S(
        \fadd_0_0_0_0_2/exponentdifferencexy [3]) );
  FADDX1 \fadd_0_0_0_0_2/sub_707/U2_4  ( .A(n5854), .B(n14553), .CI(
        \fadd_0_0_0_0_2/sub_707/carry [4]), .CO(
        \fadd_0_0_0_0_2/sub_707/carry [5]), .S(
        \fadd_0_0_0_0_2/exponentdifferencexy [4]) );
  FADDX1 \fadd_0_0_0_0_1/add_859/U1_1  ( .A(
        \fadd_0_0_0_0_1/exponentresultfar0_d2 [1]), .B(n14225), .CI(
        \fadd_0_0_0_0_1/add_859/carry [1]), .CO(
        \fadd_0_0_0_0_1/add_859/carry [2]), .S(
        \fadd_0_0_0_0_1/exponentresultfar1 [1]) );
  FADDX1 \fadd_0_0_0_0_1/add_859/U1_2  ( .A(
        \fadd_0_0_0_0_1/exponentresultfar0_d2 [2]), .B(n14225), .CI(
        \fadd_0_0_0_0_1/add_859/carry [2]), .CO(
        \fadd_0_0_0_0_1/add_859/carry [3]), .S(
        \fadd_0_0_0_0_1/exponentresultfar1 [2]) );
  FADDX1 \fadd_0_0_0_0_1/add_859/U1_3  ( .A(
        \fadd_0_0_0_0_1/exponentresultfar0_d2 [3]), .B(n14225), .CI(
        \fadd_0_0_0_0_1/add_859/carry [3]), .CO(
        \fadd_0_0_0_0_1/add_859/carry [4]), .S(
        \fadd_0_0_0_0_1/exponentresultfar1 [3]) );
  FADDX1 \fadd_0_0_0_0_1/add_859/U1_4  ( .A(
        \fadd_0_0_0_0_1/exponentresultfar0_d2 [4]), .B(n14225), .CI(
        \fadd_0_0_0_0_1/add_859/carry [4]), .CO(
        \fadd_0_0_0_0_1/add_859/carry [5]), .S(
        \fadd_0_0_0_0_1/exponentresultfar1 [4]) );
  FADDX1 \fadd_0_0_0_0_1/sub_784/U2_1  ( .A(\fadd_0_0_0_0_1/newx_d1 [5]), .B(
        n14929), .CI(\fadd_0_0_0_0_1/sub_784/carry [1]), .CO(
        \fadd_0_0_0_0_1/sub_784/carry [2]), .S(
        \fadd_0_0_0_0_1/exponentresultclose [1]) );
  FADDX1 \fadd_0_0_0_0_1/sub_784/U2_2  ( .A(\fadd_0_0_0_0_1/newx_d1 [6]), .B(
        n10411), .CI(\fadd_0_0_0_0_1/sub_784/carry [2]), .CO(
        \fadd_0_0_0_0_1/sub_784/carry [3]), .S(
        \fadd_0_0_0_0_1/exponentresultclose [2]) );
  FADDX1 \fadd_0_0_0_0_1/sub_710/U2_1  ( .A(n5911), .B(n14550), .CI(
        \fadd_0_0_0_0_1/sub_710/carry [1]), .CO(
        \fadd_0_0_0_0_1/sub_710/carry [2]), .S(
        \fadd_0_0_0_0_1/exponentdifferenceyx [1]) );
  FADDX1 \fadd_0_0_0_0_1/sub_710/U2_2  ( .A(n5912), .B(n14549), .CI(
        \fadd_0_0_0_0_1/sub_710/carry [2]), .CO(
        \fadd_0_0_0_0_1/sub_710/carry [3]), .S(
        \fadd_0_0_0_0_1/exponentdifferenceyx [2]) );
  FADDX1 \fadd_0_0_0_0_1/sub_710/U2_3  ( .A(n5913), .B(n14548), .CI(
        \fadd_0_0_0_0_1/sub_710/carry [3]), .CO(
        \fadd_0_0_0_0_1/sub_710/carry [4]), .S(
        \fadd_0_0_0_0_1/exponentdifferenceyx [3]) );
  FADDX1 \fadd_0_0_0_0_1/sub_707/U2_1  ( .A(n5923), .B(n14545), .CI(
        \fadd_0_0_0_0_1/sub_707/carry [1]), .CO(
        \fadd_0_0_0_0_1/sub_707/carry [2]), .S(
        \fadd_0_0_0_0_1/exponentdifferencexy [1]) );
  FADDX1 \fadd_0_0_0_0_1/sub_707/U2_2  ( .A(n5924), .B(n14544), .CI(
        \fadd_0_0_0_0_1/sub_707/carry [2]), .CO(
        \fadd_0_0_0_0_1/sub_707/carry [3]), .S(
        \fadd_0_0_0_0_1/exponentdifferencexy [2]) );
  FADDX1 \fadd_0_0_0_0_1/sub_707/U2_3  ( .A(n5925), .B(n14543), .CI(
        \fadd_0_0_0_0_1/sub_707/carry [3]), .CO(
        \fadd_0_0_0_0_1/sub_707/carry [4]), .S(
        \fadd_0_0_0_0_1/exponentdifferencexy [3]) );
  FADDX1 \fadd_0_0_0_0_1/sub_707/U2_4  ( .A(n5926), .B(n14542), .CI(
        \fadd_0_0_0_0_1/sub_707/carry [4]), .CO(
        \fadd_0_0_0_0_1/sub_707/carry [5]), .S(
        \fadd_0_0_0_0_1/exponentdifferencexy [4]) );
  FADDX1 \fadd_0_0_0_0_0/add_859/U1_1  ( .A(
        \fadd_0_0_0_0_0/exponentresultfar0_d2 [1]), .B(
        \fadd_0_0_0_0_0/add_859/B[1] ), .CI(\fadd_0_0_0_0_0/add_859/carry [1]), 
        .CO(\fadd_0_0_0_0_0/add_859/carry [2]), .S(
        \fadd_0_0_0_0_0/exponentresultfar1 [1]) );
  FADDX1 \fadd_0_0_0_0_0/add_859/U1_2  ( .A(
        \fadd_0_0_0_0_0/exponentresultfar0_d2 [2]), .B(
        \fadd_0_0_0_0_0/add_859/B[1] ), .CI(\fadd_0_0_0_0_0/add_859/carry [2]), 
        .CO(\fadd_0_0_0_0_0/add_859/carry [3]), .S(
        \fadd_0_0_0_0_0/exponentresultfar1 [2]) );
  FADDX1 \fadd_0_0_0_0_0/add_859/U1_3  ( .A(
        \fadd_0_0_0_0_0/exponentresultfar0_d2 [3]), .B(
        \fadd_0_0_0_0_0/add_859/B[1] ), .CI(\fadd_0_0_0_0_0/add_859/carry [3]), 
        .CO(\fadd_0_0_0_0_0/add_859/carry [4]), .S(
        \fadd_0_0_0_0_0/exponentresultfar1 [3]) );
  FADDX1 \fadd_0_0_0_0_0/add_859/U1_4  ( .A(
        \fadd_0_0_0_0_0/exponentresultfar0_d2 [4]), .B(n14224), .CI(
        \fadd_0_0_0_0_0/add_859/carry [4]), .CO(
        \fadd_0_0_0_0_0/add_859/carry [5]), .S(
        \fadd_0_0_0_0_0/exponentresultfar1 [4]) );
  FADDX1 \fadd_0_0_0_0_0/sub_784/U2_1  ( .A(\fadd_0_0_0_0_0/newx_d1 [5]), .B(
        n14928), .CI(\fadd_0_0_0_0_0/sub_784/carry [1]), .CO(
        \fadd_0_0_0_0_0/sub_784/carry [2]), .S(
        \fadd_0_0_0_0_0/exponentresultclose [1]) );
  FADDX1 \fadd_0_0_0_0_0/sub_784/U2_2  ( .A(\fadd_0_0_0_0_0/newx_d1 [6]), .B(
        n10410), .CI(\fadd_0_0_0_0_0/sub_784/carry [2]), .CO(
        \fadd_0_0_0_0_0/sub_784/carry [3]), .S(
        \fadd_0_0_0_0_0/exponentresultclose [2]) );
  FADDX1 \fadd_0_0_0_0_0/sub_710/U2_1  ( .A(n5983), .B(n14539), .CI(
        \fadd_0_0_0_0_0/sub_710/carry [1]), .CO(
        \fadd_0_0_0_0_0/sub_710/carry [2]), .S(
        \fadd_0_0_0_0_0/exponentdifferenceyx [1]) );
  FADDX1 \fadd_0_0_0_0_0/sub_710/U2_2  ( .A(n5984), .B(n14538), .CI(
        \fadd_0_0_0_0_0/sub_710/carry [2]), .CO(
        \fadd_0_0_0_0_0/sub_710/carry [3]), .S(
        \fadd_0_0_0_0_0/exponentdifferenceyx [2]) );
  FADDX1 \fadd_0_0_0_0_0/sub_710/U2_3  ( .A(n5985), .B(n14537), .CI(
        \fadd_0_0_0_0_0/sub_710/carry [3]), .CO(
        \fadd_0_0_0_0_0/sub_710/carry [4]), .S(
        \fadd_0_0_0_0_0/exponentdifferenceyx [3]) );
  FADDX1 \fadd_0_0_0_0_0/sub_707/U2_1  ( .A(n5995), .B(n14534), .CI(
        \fadd_0_0_0_0_0/sub_707/carry [1]), .CO(
        \fadd_0_0_0_0_0/sub_707/carry [2]), .S(
        \fadd_0_0_0_0_0/exponentdifferencexy [1]) );
  FADDX1 \fadd_0_0_0_0_0/sub_707/U2_2  ( .A(n5996), .B(n14533), .CI(
        \fadd_0_0_0_0_0/sub_707/carry [2]), .CO(
        \fadd_0_0_0_0_0/sub_707/carry [3]), .S(
        \fadd_0_0_0_0_0/exponentdifferencexy [2]) );
  FADDX1 \fadd_0_0_0_0_0/sub_707/U2_3  ( .A(n5997), .B(n14532), .CI(
        \fadd_0_0_0_0_0/sub_707/carry [3]), .CO(
        \fadd_0_0_0_0_0/sub_707/carry [4]), .S(
        \fadd_0_0_0_0_0/exponentdifferencexy [3]) );
  FADDX1 \fadd_0_0_0_0_0/sub_707/U2_4  ( .A(n5998), .B(n14531), .CI(
        \fadd_0_0_0_0_0/sub_707/carry [4]), .CO(
        \fadd_0_0_0_0_0/sub_707/carry [5]), .S(
        \fadd_0_0_0_0_0/exponentdifferencexy [4]) );
  FADDX1 \add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/U1_1  ( .A(
        \add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/A[1] ), .B(
        \add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/B[1] ), .CI(
        \add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/carry [1]), .CO(
        \add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/carry [2]), .S(
        \fmul_0_0_0_0_0/exppostnorm [1]) );
  FADDX1 \add_2_root_sub_1_root_fmul_0_0_0_0_0/add_321/U1_1  ( .A(n5959), .B(
        n5947), .CI(\add_2_root_sub_1_root_fmul_0_0_0_0_0/add_321/carry [1]), 
        .CO(\add_2_root_sub_1_root_fmul_0_0_0_0_0/add_321/carry [2]), .S(
        \add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/A[1] ) );
  FADDX1 \add_2_root_sub_1_root_fmul_0_0_0_0_0/add_321/U1_2  ( .A(n5960), .B(
        n5948), .CI(\add_2_root_sub_1_root_fmul_0_0_0_0_0/add_321/carry [2]), 
        .CO(\add_2_root_sub_1_root_fmul_0_0_0_0_0/add_321/carry [3]), .S(
        \add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/A[2] ) );
  FADDX1 \add_2_root_sub_1_root_fmul_0_0_0_0_0/add_321/U1_3  ( .A(n5961), .B(
        n5949), .CI(\add_2_root_sub_1_root_fmul_0_0_0_0_0/add_321/carry [3]), 
        .CO(\add_2_root_sub_1_root_fmul_0_0_0_0_0/add_321/carry [4]), .S(
        \add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/A[3] ) );
  FADDX1 \add_2_root_sub_1_root_fmul_0_0_0_0_0/add_321/U1_4  ( .A(n5962), .B(
        n5950), .CI(\add_2_root_sub_1_root_fmul_0_0_0_0_0/add_321/carry [4]), 
        .CO(\add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/A[5] ), .S(
        \add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/A[4] ) );
  FADDX1 \add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/U1_1  ( .A(
        \add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/A[1] ), .B(
        \add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/B[1] ), .CI(
        \add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/carry [1]), .CO(
        \add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/carry [2]), .S(
        \fmul_0_0_0_0_1/exppostnorm [1]) );
  FADDX1 \add_2_root_sub_1_root_fmul_0_0_0_0_1/add_321/U1_1  ( .A(n5887), .B(
        n5875), .CI(\add_2_root_sub_1_root_fmul_0_0_0_0_1/add_321/carry [1]), 
        .CO(\add_2_root_sub_1_root_fmul_0_0_0_0_1/add_321/carry [2]), .S(
        \add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/A[1] ) );
  FADDX1 \add_2_root_sub_1_root_fmul_0_0_0_0_1/add_321/U1_2  ( .A(n5888), .B(
        n5876), .CI(\add_2_root_sub_1_root_fmul_0_0_0_0_1/add_321/carry [2]), 
        .CO(\add_2_root_sub_1_root_fmul_0_0_0_0_1/add_321/carry [3]), .S(
        \add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/A[2] ) );
  FADDX1 \add_2_root_sub_1_root_fmul_0_0_0_0_1/add_321/U1_3  ( .A(n5889), .B(
        n5877), .CI(\add_2_root_sub_1_root_fmul_0_0_0_0_1/add_321/carry [3]), 
        .CO(\add_2_root_sub_1_root_fmul_0_0_0_0_1/add_321/carry [4]), .S(
        \add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/A[3] ) );
  FADDX1 \add_2_root_sub_1_root_fmul_0_0_0_0_1/add_321/U1_4  ( .A(n5890), .B(
        n5878), .CI(\add_2_root_sub_1_root_fmul_0_0_0_0_1/add_321/carry [4]), 
        .CO(\add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/A[5] ), .S(
        \add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/A[4] ) );
  FADDX1 \add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/U1_1  ( .A(
        \add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/A[1] ), .B(
        \add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/B[1] ), .CI(
        \add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/carry [1]), .CO(
        \add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/carry [2]), .S(
        \fmul_0_0_0_0_2/exppostnorm [1]) );
  FADDX1 \add_2_root_sub_1_root_fmul_0_0_0_0_2/add_321/U1_1  ( .A(n5815), .B(
        n5803), .CI(\add_2_root_sub_1_root_fmul_0_0_0_0_2/add_321/carry [1]), 
        .CO(\add_2_root_sub_1_root_fmul_0_0_0_0_2/add_321/carry [2]), .S(
        \add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/A[1] ) );
  FADDX1 \add_2_root_sub_1_root_fmul_0_0_0_0_2/add_321/U1_2  ( .A(n5816), .B(
        n5804), .CI(\add_2_root_sub_1_root_fmul_0_0_0_0_2/add_321/carry [2]), 
        .CO(\add_2_root_sub_1_root_fmul_0_0_0_0_2/add_321/carry [3]), .S(
        \add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/A[2] ) );
  FADDX1 \add_2_root_sub_1_root_fmul_0_0_0_0_2/add_321/U1_3  ( .A(n5817), .B(
        n5805), .CI(\add_2_root_sub_1_root_fmul_0_0_0_0_2/add_321/carry [3]), 
        .CO(\add_2_root_sub_1_root_fmul_0_0_0_0_2/add_321/carry [4]), .S(
        \add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/A[3] ) );
  FADDX1 \add_2_root_sub_1_root_fmul_0_0_0_0_2/add_321/U1_4  ( .A(n5818), .B(
        n5806), .CI(\add_2_root_sub_1_root_fmul_0_0_0_0_2/add_321/carry [4]), 
        .CO(\add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/A[5] ), .S(
        \add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/A[4] ) );
  FADDX1 \add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/U1_1  ( .A(
        \add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/A[1] ), .B(
        \add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/B[1] ), .CI(
        \add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/carry [1]), .CO(
        \add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/carry [2]), .S(
        \fmul_0_0_0_0_3/exppostnorm [1]) );
  FADDX1 \add_2_root_sub_1_root_fmul_0_0_0_0_3/add_321/U1_1  ( .A(n5743), .B(
        n5731), .CI(\add_2_root_sub_1_root_fmul_0_0_0_0_3/add_321/carry [1]), 
        .CO(\add_2_root_sub_1_root_fmul_0_0_0_0_3/add_321/carry [2]), .S(
        \add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/A[1] ) );
  FADDX1 \add_2_root_sub_1_root_fmul_0_0_0_0_3/add_321/U1_2  ( .A(n5744), .B(
        n5732), .CI(\add_2_root_sub_1_root_fmul_0_0_0_0_3/add_321/carry [2]), 
        .CO(\add_2_root_sub_1_root_fmul_0_0_0_0_3/add_321/carry [3]), .S(
        \add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/A[2] ) );
  FADDX1 \add_2_root_sub_1_root_fmul_0_0_0_0_3/add_321/U1_3  ( .A(n5745), .B(
        n5733), .CI(\add_2_root_sub_1_root_fmul_0_0_0_0_3/add_321/carry [3]), 
        .CO(\add_2_root_sub_1_root_fmul_0_0_0_0_3/add_321/carry [4]), .S(
        \add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/A[3] ) );
  FADDX1 \add_2_root_sub_1_root_fmul_0_0_0_0_3/add_321/U1_4  ( .A(n5746), .B(
        n5734), .CI(\add_2_root_sub_1_root_fmul_0_0_0_0_3/add_321/carry [4]), 
        .CO(\add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/A[5] ), .S(
        \add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/A[4] ) );
  FADDX1 \add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/U1_1  ( .A(
        \add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/A[1] ), .B(
        \add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/B[1] ), .CI(
        \add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/carry [1]), .CO(
        \add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/carry [2]), .S(
        \fmul_0_0_0_0_4/exppostnorm [1]) );
  FADDX1 \add_2_root_sub_1_root_fmul_0_0_0_0_4/add_321/U1_1  ( .A(n5671), .B(
        n5659), .CI(\add_2_root_sub_1_root_fmul_0_0_0_0_4/add_321/carry [1]), 
        .CO(\add_2_root_sub_1_root_fmul_0_0_0_0_4/add_321/carry [2]), .S(
        \add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/A[1] ) );
  FADDX1 \add_2_root_sub_1_root_fmul_0_0_0_0_4/add_321/U1_2  ( .A(n5672), .B(
        n5660), .CI(\add_2_root_sub_1_root_fmul_0_0_0_0_4/add_321/carry [2]), 
        .CO(\add_2_root_sub_1_root_fmul_0_0_0_0_4/add_321/carry [3]), .S(
        \add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/A[2] ) );
  FADDX1 \add_2_root_sub_1_root_fmul_0_0_0_0_4/add_321/U1_3  ( .A(n5673), .B(
        n5661), .CI(\add_2_root_sub_1_root_fmul_0_0_0_0_4/add_321/carry [3]), 
        .CO(\add_2_root_sub_1_root_fmul_0_0_0_0_4/add_321/carry [4]), .S(
        \add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/A[3] ) );
  FADDX1 \add_2_root_sub_1_root_fmul_0_0_0_0_4/add_321/U1_4  ( .A(n5674), .B(
        n5662), .CI(\add_2_root_sub_1_root_fmul_0_0_0_0_4/add_321/carry [4]), 
        .CO(\add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/A[5] ), .S(
        \add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/A[4] ) );
  FADDX1 \add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/U1_1  ( .A(
        \add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/A[1] ), .B(
        \add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/B[1] ), .CI(
        \add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/carry [1]), .CO(
        \add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/carry [2]), .S(
        \fmul_0_0_0_0_5/exppostnorm [1]) );
  FADDX1 \add_2_root_sub_1_root_fmul_0_0_0_0_5/add_321/U1_1  ( .A(n5599), .B(
        n5587), .CI(\add_2_root_sub_1_root_fmul_0_0_0_0_5/add_321/carry [1]), 
        .CO(\add_2_root_sub_1_root_fmul_0_0_0_0_5/add_321/carry [2]), .S(
        \add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/A[1] ) );
  FADDX1 \add_2_root_sub_1_root_fmul_0_0_0_0_5/add_321/U1_2  ( .A(n5600), .B(
        n5588), .CI(\add_2_root_sub_1_root_fmul_0_0_0_0_5/add_321/carry [2]), 
        .CO(\add_2_root_sub_1_root_fmul_0_0_0_0_5/add_321/carry [3]), .S(
        \add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/A[2] ) );
  FADDX1 \add_2_root_sub_1_root_fmul_0_0_0_0_5/add_321/U1_3  ( .A(n5601), .B(
        n5589), .CI(\add_2_root_sub_1_root_fmul_0_0_0_0_5/add_321/carry [3]), 
        .CO(\add_2_root_sub_1_root_fmul_0_0_0_0_5/add_321/carry [4]), .S(
        \add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/A[3] ) );
  FADDX1 \add_2_root_sub_1_root_fmul_0_0_0_0_5/add_321/U1_4  ( .A(n5602), .B(
        n5590), .CI(\add_2_root_sub_1_root_fmul_0_0_0_0_5/add_321/carry [4]), 
        .CO(\add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/A[5] ), .S(
        \add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/A[4] ) );
  FADDX1 \add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/U1_1  ( .A(
        \add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/A[1] ), .B(
        \add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/B[1] ), .CI(
        \add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/carry [1]), .CO(
        \add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/carry [2]), .S(
        \fmul_0_0_0_0_6/exppostnorm [1]) );
  FADDX1 \add_2_root_sub_1_root_fmul_0_0_0_0_6/add_321/U1_1  ( .A(n5527), .B(
        n5515), .CI(\add_2_root_sub_1_root_fmul_0_0_0_0_6/add_321/carry [1]), 
        .CO(\add_2_root_sub_1_root_fmul_0_0_0_0_6/add_321/carry [2]), .S(
        \add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/A[1] ) );
  FADDX1 \add_2_root_sub_1_root_fmul_0_0_0_0_6/add_321/U1_2  ( .A(n5528), .B(
        n5516), .CI(\add_2_root_sub_1_root_fmul_0_0_0_0_6/add_321/carry [2]), 
        .CO(\add_2_root_sub_1_root_fmul_0_0_0_0_6/add_321/carry [3]), .S(
        \add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/A[2] ) );
  FADDX1 \add_2_root_sub_1_root_fmul_0_0_0_0_6/add_321/U1_3  ( .A(n5529), .B(
        n5517), .CI(\add_2_root_sub_1_root_fmul_0_0_0_0_6/add_321/carry [3]), 
        .CO(\add_2_root_sub_1_root_fmul_0_0_0_0_6/add_321/carry [4]), .S(
        \add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/A[3] ) );
  FADDX1 \add_2_root_sub_1_root_fmul_0_0_0_0_6/add_321/U1_4  ( .A(n5530), .B(
        n5518), .CI(\add_2_root_sub_1_root_fmul_0_0_0_0_6/add_321/carry [4]), 
        .CO(\add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/A[5] ), .S(
        \add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/A[4] ) );
  FADDX1 \add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/U1_1  ( .A(
        \add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/A[1] ), .B(
        \add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/B[1] ), .CI(
        \add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/carry [1]), .CO(
        \add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/carry [2]), .S(
        \fmul_0_0_0_0_7/exppostnorm [1]) );
  FADDX1 \add_2_root_sub_1_root_fmul_0_0_0_0_7/add_321/U1_1  ( .A(n5455), .B(
        n5443), .CI(\add_2_root_sub_1_root_fmul_0_0_0_0_7/add_321/carry [1]), 
        .CO(\add_2_root_sub_1_root_fmul_0_0_0_0_7/add_321/carry [2]), .S(
        \add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/A[1] ) );
  FADDX1 \add_2_root_sub_1_root_fmul_0_0_0_0_7/add_321/U1_2  ( .A(n5456), .B(
        n5444), .CI(\add_2_root_sub_1_root_fmul_0_0_0_0_7/add_321/carry [2]), 
        .CO(\add_2_root_sub_1_root_fmul_0_0_0_0_7/add_321/carry [3]), .S(
        \add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/A[2] ) );
  FADDX1 \add_2_root_sub_1_root_fmul_0_0_0_0_7/add_321/U1_3  ( .A(n5457), .B(
        n5445), .CI(\add_2_root_sub_1_root_fmul_0_0_0_0_7/add_321/carry [3]), 
        .CO(\add_2_root_sub_1_root_fmul_0_0_0_0_7/add_321/carry [4]), .S(
        \add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/A[3] ) );
  FADDX1 \add_2_root_sub_1_root_fmul_0_0_0_0_7/add_321/U1_4  ( .A(n5458), .B(
        n5446), .CI(\add_2_root_sub_1_root_fmul_0_0_0_0_7/add_321/carry [4]), 
        .CO(\add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/A[5] ), .S(
        \add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/A[4] ) );
  FADDX1 \add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/U1_1  ( .A(
        \add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/A[1] ), .B(
        \add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/B[1] ), .CI(
        \add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/carry [1]), .CO(
        \add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/carry [2]), .S(
        \fmul_0_0_0_0_8/exppostnorm [1]) );
  FADDX1 \add_2_root_sub_1_root_fmul_0_0_0_0_8/add_321/U1_1  ( .A(n5383), .B(
        n5371), .CI(\add_2_root_sub_1_root_fmul_0_0_0_0_8/add_321/carry [1]), 
        .CO(\add_2_root_sub_1_root_fmul_0_0_0_0_8/add_321/carry [2]), .S(
        \add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/A[1] ) );
  FADDX1 \add_2_root_sub_1_root_fmul_0_0_0_0_8/add_321/U1_2  ( .A(n5384), .B(
        n5372), .CI(\add_2_root_sub_1_root_fmul_0_0_0_0_8/add_321/carry [2]), 
        .CO(\add_2_root_sub_1_root_fmul_0_0_0_0_8/add_321/carry [3]), .S(
        \add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/A[2] ) );
  FADDX1 \add_2_root_sub_1_root_fmul_0_0_0_0_8/add_321/U1_3  ( .A(n5385), .B(
        n5373), .CI(\add_2_root_sub_1_root_fmul_0_0_0_0_8/add_321/carry [3]), 
        .CO(\add_2_root_sub_1_root_fmul_0_0_0_0_8/add_321/carry [4]), .S(
        \add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/A[3] ) );
  FADDX1 \add_2_root_sub_1_root_fmul_0_0_0_0_8/add_321/U1_4  ( .A(n5386), .B(
        n5374), .CI(\add_2_root_sub_1_root_fmul_0_0_0_0_8/add_321/carry [4]), 
        .CO(\add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/A[5] ), .S(
        \add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/A[4] ) );
  FADDX1 \add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/U1_1  ( .A(
        \add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/A[1] ), .B(
        \add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/B[1] ), .CI(
        \add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/carry [1]), .CO(
        \add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/carry [2]), .S(
        \fmul_0_0_0_0_9/exppostnorm [1]) );
  FADDX1 \add_2_root_sub_1_root_fmul_0_0_0_0_9/add_321/U1_1  ( .A(n5311), .B(
        n5299), .CI(\add_2_root_sub_1_root_fmul_0_0_0_0_9/add_321/carry [1]), 
        .CO(\add_2_root_sub_1_root_fmul_0_0_0_0_9/add_321/carry [2]), .S(
        \add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/A[1] ) );
  FADDX1 \add_2_root_sub_1_root_fmul_0_0_0_0_9/add_321/U1_2  ( .A(n5312), .B(
        n5300), .CI(\add_2_root_sub_1_root_fmul_0_0_0_0_9/add_321/carry [2]), 
        .CO(\add_2_root_sub_1_root_fmul_0_0_0_0_9/add_321/carry [3]), .S(
        \add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/A[2] ) );
  FADDX1 \add_2_root_sub_1_root_fmul_0_0_0_0_9/add_321/U1_3  ( .A(n5313), .B(
        n5301), .CI(\add_2_root_sub_1_root_fmul_0_0_0_0_9/add_321/carry [3]), 
        .CO(\add_2_root_sub_1_root_fmul_0_0_0_0_9/add_321/carry [4]), .S(
        \add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/A[3] ) );
  FADDX1 \add_2_root_sub_1_root_fmul_0_0_0_0_9/add_321/U1_4  ( .A(n5314), .B(
        n5302), .CI(\add_2_root_sub_1_root_fmul_0_0_0_0_9/add_321/carry [4]), 
        .CO(\add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/A[5] ), .S(
        \add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/A[4] ) );
  FADDX1 \sub_0_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_300/U2_1  ( 
        .A(
        \add_0_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .B(n14527), .CI(n14526), .CO(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [2]), .S(\fadd_0_0_0_0_8/fracrclosexmy [1]) );
  FADDX1 \sub_0_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_300/U2_3  ( 
        .A(\fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ), .B(
        n14530), .CI(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [3]), .CO(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [4]), .S(\fadd_0_0_0_0_8/fracrclosexmy [3]) );
  FADDX1 \sub_0_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_300/U2_4  ( 
        .A(\fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ), .B(
        n14529), .CI(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [4]), .CO(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [5]), .S(\fadd_0_0_0_0_8/fracrclosexmy [4]) );
  FADDX1 \add_0_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_303/U1_2  ( 
        .A(\fadd_0_0_0_0_8/fracyclose1 [2]), .B(
        \add_0_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[2] ), .CI(
        \add_0_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [2]), .CO(
        \add_0_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [3]), .S(\fadd_0_0_0_0_8/fracrcloseymx [2]) );
  FADDX1 \add_0_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_303/U1_3  ( 
        .A(\fadd_0_0_0_0_8/fracyclose1 [3]), .B(
        \add_0_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[3] ), .CI(
        \add_0_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [3]), .CO(
        \add_0_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [4]), .S(\fadd_0_0_0_0_8/fracrcloseymx [3]) );
  FADDX1 \add_0_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_303/U1_4  ( 
        .A(\fadd_0_0_0_0_8/fracyclose1 [4]), .B(
        \add_0_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[4] ), .CI(
        \add_0_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [4]), .CO(
        \add_0_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [5]), .S(\fadd_0_0_0_0_8/fracrcloseymx [4]) );
  FADDX1 \sub_0_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_300/U2_1  ( 
        .A(
        \add_0_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .B(n14518), .CI(n14517), .CO(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [2]), .S(\fadd_0_0_0_0_9/fracrclosexmy [1]) );
  FADDX1 \sub_0_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_300/U2_3  ( 
        .A(\fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ), .B(
        n14521), .CI(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [3]), .CO(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [4]), .S(\fadd_0_0_0_0_9/fracrclosexmy [3]) );
  FADDX1 \sub_0_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_300/U2_4  ( 
        .A(\fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ), .B(
        n14520), .CI(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [4]), .CO(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [5]), .S(\fadd_0_0_0_0_9/fracrclosexmy [4]) );
  FADDX1 \add_0_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_303/U1_2  ( 
        .A(\fadd_0_0_0_0_9/fracyclose1 [2]), .B(
        \add_0_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[2] ), .CI(
        \add_0_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [2]), .CO(
        \add_0_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [3]), .S(\fadd_0_0_0_0_9/fracrcloseymx [2]) );
  FADDX1 \add_0_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_303/U1_3  ( 
        .A(\fadd_0_0_0_0_9/fracyclose1 [3]), .B(
        \add_0_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[3] ), .CI(
        \add_0_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [3]), .CO(
        \add_0_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [4]), .S(\fadd_0_0_0_0_9/fracrcloseymx [3]) );
  FADDX1 \add_0_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_303/U1_4  ( 
        .A(\fadd_0_0_0_0_9/fracyclose1 [4]), .B(
        \add_0_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[4] ), .CI(
        \add_0_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [4]), .CO(
        \add_0_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [5]), .S(\fadd_0_0_0_0_9/fracrcloseymx [4]) );
  FADDX1 \sub_0_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_300/U2_1  ( 
        .A(
        \add_0_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .B(n14509), .CI(n14508), .CO(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [2]), .S(\fadd_0_0_0_0_0/fracrclosexmy [1]) );
  FADDX1 \sub_0_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_300/U2_2  ( 
        .A(\fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ), .B(
        n14510), .CI(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [2]), .CO(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [3]), .S(\fadd_0_0_0_0_0/fracrclosexmy [2]) );
  FADDX1 \sub_0_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_300/U2_3  ( 
        .A(\fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ), .B(
        n14512), .CI(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [3]), .CO(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [4]), .S(\fadd_0_0_0_0_0/fracrclosexmy [3]) );
  FADDX1 \sub_0_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_300/U2_4  ( 
        .A(\fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ), .B(
        n14511), .CI(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [4]), .CO(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [5]), .S(\fadd_0_0_0_0_0/fracrclosexmy [4]) );
  FADDX1 \add_0_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_303/U1_2  ( 
        .A(\fadd_0_0_0_0_0/fracyclose1 [2]), .B(
        \add_0_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[2] ), .CI(
        \add_0_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [2]), .CO(
        \add_0_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [3]), .S(\fadd_0_0_0_0_0/fracrcloseymx [2]) );
  FADDX1 \add_0_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_303/U1_3  ( 
        .A(\fadd_0_0_0_0_0/fracyclose1 [3]), .B(
        \add_0_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[3] ), .CI(
        \add_0_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [3]), .CO(
        \add_0_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [4]), .S(\fadd_0_0_0_0_0/fracrcloseymx [3]) );
  FADDX1 \add_0_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_303/U1_4  ( 
        .A(\fadd_0_0_0_0_0/fracyclose1 [4]), .B(
        \add_0_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[4] ), .CI(
        \add_0_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [4]), .CO(
        \add_0_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [5]), .S(\fadd_0_0_0_0_0/fracrcloseymx [4]) );
  FADDX1 \sub_0_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_300/U2_1  ( 
        .A(
        \add_0_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .B(n14500), .CI(n14499), .CO(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [2]), .S(\fadd_0_0_0_0_4/fracrclosexmy [1]) );
  FADDX1 \sub_0_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_300/U2_2  ( 
        .A(\fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ), .B(
        n14501), .CI(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [2]), .CO(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [3]), .S(\fadd_0_0_0_0_4/fracrclosexmy [2]) );
  FADDX1 \sub_0_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_300/U2_3  ( 
        .A(\fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ), .B(
        n14503), .CI(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [3]), .CO(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [4]), .S(\fadd_0_0_0_0_4/fracrclosexmy [3]) );
  FADDX1 \sub_0_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_300/U2_4  ( 
        .A(\fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ), .B(
        n14502), .CI(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [4]), .CO(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [5]), .S(\fadd_0_0_0_0_4/fracrclosexmy [4]) );
  FADDX1 \add_0_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_303/U1_2  ( 
        .A(\fadd_0_0_0_0_4/fracyclose1 [2]), .B(
        \add_0_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[2] ), .CI(
        \add_0_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [2]), .CO(
        \add_0_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [3]), .S(\fadd_0_0_0_0_4/fracrcloseymx [2]) );
  FADDX1 \add_0_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_303/U1_3  ( 
        .A(\fadd_0_0_0_0_4/fracyclose1 [3]), .B(
        \add_0_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[3] ), .CI(
        \add_0_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [3]), .CO(
        \add_0_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [4]), .S(\fadd_0_0_0_0_4/fracrcloseymx [3]) );
  FADDX1 \add_0_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_303/U1_4  ( 
        .A(\fadd_0_0_0_0_4/fracyclose1 [4]), .B(
        \add_0_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[4] ), .CI(
        \add_0_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [4]), .CO(
        \add_0_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [5]), .S(\fadd_0_0_0_0_4/fracrcloseymx [4]) );
  FADDX1 \sub_0_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_300/U2_1  ( 
        .A(
        \add_0_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .B(n14491), .CI(n14490), .CO(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [2]), .S(\fadd_0_0_0_0_6/fracrclosexmy [1]) );
  FADDX1 \sub_0_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_300/U2_3  ( 
        .A(\fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ), .B(
        n14494), .CI(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [3]), .CO(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [4]), .S(\fadd_0_0_0_0_6/fracrclosexmy [3]) );
  FADDX1 \sub_0_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_300/U2_4  ( 
        .A(\fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ), .B(
        n14493), .CI(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [4]), .CO(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [5]), .S(\fadd_0_0_0_0_6/fracrclosexmy [4]) );
  FADDX1 \add_0_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_303/U1_2  ( 
        .A(\fadd_0_0_0_0_6/fracyclose1 [2]), .B(
        \add_0_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[2] ), .CI(
        \add_0_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [2]), .CO(
        \add_0_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [3]), .S(\fadd_0_0_0_0_6/fracrcloseymx [2]) );
  FADDX1 \add_0_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_303/U1_3  ( 
        .A(\fadd_0_0_0_0_6/fracyclose1 [3]), .B(
        \add_0_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[3] ), .CI(
        \add_0_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [3]), .CO(
        \add_0_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [4]), .S(\fadd_0_0_0_0_6/fracrcloseymx [3]) );
  FADDX1 \add_0_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_303/U1_4  ( 
        .A(\fadd_0_0_0_0_6/fracyclose1 [4]), .B(
        \add_0_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[4] ), .CI(
        \add_0_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [4]), .CO(
        \add_0_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [5]), .S(\fadd_0_0_0_0_6/fracrcloseymx [4]) );
  FADDX1 \sub_0_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_300/U2_1  ( 
        .A(
        \add_0_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .B(n14482), .CI(n14481), .CO(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [2]), .S(\fadd_0_0_0_0_7/fracrclosexmy [1]) );
  FADDX1 \sub_0_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_300/U2_3  ( 
        .A(\fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ), .B(
        n14485), .CI(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [3]), .CO(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [4]), .S(\fadd_0_0_0_0_7/fracrclosexmy [3]) );
  FADDX1 \sub_0_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_300/U2_4  ( 
        .A(\fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ), .B(
        n14484), .CI(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [4]), .CO(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [5]), .S(\fadd_0_0_0_0_7/fracrclosexmy [4]) );
  FADDX1 \add_0_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_303/U1_2  ( 
        .A(\fadd_0_0_0_0_7/fracyclose1 [2]), .B(
        \add_0_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[2] ), .CI(
        \add_0_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [2]), .CO(
        \add_0_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [3]), .S(\fadd_0_0_0_0_7/fracrcloseymx [2]) );
  FADDX1 \add_0_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_303/U1_3  ( 
        .A(\fadd_0_0_0_0_7/fracyclose1 [3]), .B(
        \add_0_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[3] ), .CI(
        \add_0_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [3]), .CO(
        \add_0_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [4]), .S(\fadd_0_0_0_0_7/fracrcloseymx [3]) );
  FADDX1 \add_0_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_303/U1_4  ( 
        .A(\fadd_0_0_0_0_7/fracyclose1 [4]), .B(
        \add_0_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[4] ), .CI(
        \add_0_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [4]), .CO(
        \add_0_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [5]), .S(\fadd_0_0_0_0_7/fracrcloseymx [4]) );
  FADDX1 \sub_0_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_300/U2_1  ( 
        .A(
        \add_0_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .B(n14473), .CI(n14472), .CO(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [2]), .S(\fadd_0_0_0_0_5/fracrclosexmy [1]) );
  FADDX1 \sub_0_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_300/U2_2  ( 
        .A(\fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ), .B(
        n14474), .CI(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [2]), .CO(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [3]), .S(\fadd_0_0_0_0_5/fracrclosexmy [2]) );
  FADDX1 \sub_0_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_300/U2_3  ( 
        .A(\fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ), .B(
        n14476), .CI(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [3]), .CO(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [4]), .S(\fadd_0_0_0_0_5/fracrclosexmy [3]) );
  FADDX1 \sub_0_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_300/U2_4  ( 
        .A(\fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ), .B(
        n14475), .CI(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [4]), .CO(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [5]), .S(\fadd_0_0_0_0_5/fracrclosexmy [4]) );
  FADDX1 \add_0_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_303/U1_2  ( 
        .A(\fadd_0_0_0_0_5/fracyclose1 [2]), .B(
        \add_0_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[2] ), .CI(
        \add_0_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [2]), .CO(
        \add_0_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [3]), .S(\fadd_0_0_0_0_5/fracrcloseymx [2]) );
  FADDX1 \add_0_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_303/U1_3  ( 
        .A(\fadd_0_0_0_0_5/fracyclose1 [3]), .B(
        \add_0_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[3] ), .CI(
        \add_0_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [3]), .CO(
        \add_0_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [4]), .S(\fadd_0_0_0_0_5/fracrcloseymx [3]) );
  FADDX1 \add_0_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_303/U1_4  ( 
        .A(\fadd_0_0_0_0_5/fracyclose1 [4]), .B(
        \add_0_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[4] ), .CI(
        \add_0_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [4]), .CO(
        \add_0_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [5]), .S(\fadd_0_0_0_0_5/fracrcloseymx [4]) );
  FADDX1 \sub_0_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_300/U2_1  ( 
        .A(
        \add_0_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .B(n14464), .CI(n14463), .CO(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [2]), .S(\fadd_0_0_0_0_2/fracrclosexmy [1]) );
  FADDX1 \sub_0_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_300/U2_2  ( 
        .A(\fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ), .B(
        n14465), .CI(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [2]), .CO(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [3]), .S(\fadd_0_0_0_0_2/fracrclosexmy [2]) );
  FADDX1 \sub_0_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_300/U2_3  ( 
        .A(\fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ), .B(
        n14467), .CI(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [3]), .CO(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [4]), .S(\fadd_0_0_0_0_2/fracrclosexmy [3]) );
  FADDX1 \sub_0_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_300/U2_4  ( 
        .A(\fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ), .B(
        n14466), .CI(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [4]), .CO(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [5]), .S(\fadd_0_0_0_0_2/fracrclosexmy [4]) );
  FADDX1 \add_0_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_303/U1_2  ( 
        .A(\fadd_0_0_0_0_2/fracyclose1 [2]), .B(
        \add_0_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[2] ), .CI(
        \add_0_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [2]), .CO(
        \add_0_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [3]), .S(\fadd_0_0_0_0_2/fracrcloseymx [2]) );
  FADDX1 \add_0_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_303/U1_3  ( 
        .A(\fadd_0_0_0_0_2/fracyclose1 [3]), .B(
        \add_0_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[3] ), .CI(
        \add_0_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [3]), .CO(
        \add_0_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [4]), .S(\fadd_0_0_0_0_2/fracrcloseymx [3]) );
  FADDX1 \add_0_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_303/U1_4  ( 
        .A(\fadd_0_0_0_0_2/fracyclose1 [4]), .B(
        \add_0_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[4] ), .CI(
        \add_0_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [4]), .CO(
        \add_0_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [5]), .S(\fadd_0_0_0_0_2/fracrcloseymx [4]) );
  FADDX1 \sub_0_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_300/U2_1  ( 
        .A(
        \add_0_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .B(n14455), .CI(n14454), .CO(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [2]), .S(\fadd_0_0_0_0_3/fracrclosexmy [1]) );
  FADDX1 \sub_0_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_300/U2_3  ( 
        .A(\fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ), .B(
        n14458), .CI(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [3]), .CO(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [4]), .S(\fadd_0_0_0_0_3/fracrclosexmy [3]) );
  FADDX1 \sub_0_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_300/U2_4  ( 
        .A(\fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ), .B(
        n14457), .CI(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [4]), .CO(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [5]), .S(\fadd_0_0_0_0_3/fracrclosexmy [4]) );
  FADDX1 \add_0_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_303/U1_2  ( 
        .A(\fadd_0_0_0_0_3/fracyclose1 [2]), .B(
        \add_0_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[2] ), .CI(
        \add_0_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [2]), .CO(
        \add_0_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [3]), .S(\fadd_0_0_0_0_3/fracrcloseymx [2]) );
  FADDX1 \add_0_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_303/U1_3  ( 
        .A(\fadd_0_0_0_0_3/fracyclose1 [3]), .B(
        \add_0_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[3] ), .CI(
        \add_0_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [3]), .CO(
        \add_0_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [4]), .S(\fadd_0_0_0_0_3/fracrcloseymx [3]) );
  FADDX1 \add_0_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_303/U1_4  ( 
        .A(\fadd_0_0_0_0_3/fracyclose1 [4]), .B(
        \add_0_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[4] ), .CI(
        \add_0_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [4]), .CO(
        \add_0_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [5]), .S(\fadd_0_0_0_0_3/fracrcloseymx [4]) );
  FADDX1 \sub_0_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_300/U2_1  ( 
        .A(
        \add_0_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .B(n14446), .CI(n14445), .CO(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [2]), .S(\fadd_0_0_0_0_1/fracrclosexmy [1]) );
  FADDX1 \sub_0_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_300/U2_2  ( 
        .A(\fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ), .B(
        n14447), .CI(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [2]), .CO(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [3]), .S(\fadd_0_0_0_0_1/fracrclosexmy [2]) );
  FADDX1 \sub_0_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_300/U2_3  ( 
        .A(\fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ), .B(
        n14449), .CI(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [3]), .CO(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [4]), .S(\fadd_0_0_0_0_1/fracrclosexmy [3]) );
  FADDX1 \sub_0_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_300/U2_4  ( 
        .A(\fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ), .B(
        n14448), .CI(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [4]), .CO(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [5]), .S(\fadd_0_0_0_0_1/fracrclosexmy [4]) );
  FADDX1 \add_0_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_303/U1_2  ( 
        .A(\fadd_0_0_0_0_1/fracyclose1 [2]), .B(
        \add_0_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[2] ), .CI(
        \add_0_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [2]), .CO(
        \add_0_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [3]), .S(\fadd_0_0_0_0_1/fracrcloseymx [2]) );
  FADDX1 \add_0_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_303/U1_3  ( 
        .A(\fadd_0_0_0_0_1/fracyclose1 [3]), .B(
        \add_0_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[3] ), .CI(
        \add_0_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [3]), .CO(
        \add_0_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [4]), .S(\fadd_0_0_0_0_1/fracrcloseymx [3]) );
  FADDX1 \add_0_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_303/U1_4  ( 
        .A(\fadd_0_0_0_0_1/fracyclose1 [4]), .B(
        \add_0_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[4] ), .CI(
        \add_0_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [4]), .CO(
        \add_0_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [5]), .S(\fadd_0_0_0_0_1/fracrcloseymx [4]) );
  DFFX1 \current_fsm_reg[53]  ( .D(\U4/Z_53 ), .CLK(clk), .Q(n13748), .QN(
        n12007) );
  DFFX1 \current_fsm_reg[49]  ( .D(\U4/Z_49 ), .CLK(clk), .Q(n13587), .QN(
        n12143) );
  DFFX1 \current_fsm_reg[48]  ( .D(\U4/Z_48 ), .CLK(clk), .Q(n13586), .QN(
        n12009) );
  DFFX1 \current_fsm_reg[50]  ( .D(\U4/Z_50 ), .CLK(clk), .Q(n13497), .QN(
        n11959) );
  DFFX1 \fadd_0_0_0_0_1/n279_q_reg  ( .D(\fadd_0_0_0_0_1/selectclosepath_d1 ), 
        .CLK(clk), .Q(n13649), .QN(n12839) );
  DFFX1 \fadd_0_0_0_0_3/n279_q_reg  ( .D(\fadd_0_0_0_0_3/selectclosepath_d1 ), 
        .CLK(clk), .Q(n13650), .QN(n12841) );
  DFFX1 \fadd_0_0_0_0_9/n279_q_reg  ( .D(\fadd_0_0_0_0_9/selectclosepath_d1 ), 
        .CLK(clk), .Q(n13653), .QN(n12847) );
  DFFX1 \fadd_0_0_0_0_5/n279_q_reg  ( .D(\fadd_0_0_0_0_5/selectclosepath_d1 ), 
        .CLK(clk), .Q(n13651), .QN(n12843) );
  DFFX1 \fadd_0_0_0_0_7/n279_q_reg  ( .D(\fadd_0_0_0_0_7/selectclosepath_d1 ), 
        .CLK(clk), .Q(n13652), .QN(n12845) );
  DFFX1 \fadd_0_0_0_0_6/n279_q_reg  ( .D(\fadd_0_0_0_0_6/selectclosepath_d1 ), 
        .CLK(clk), .Q(n13647), .QN(n12844) );
  DFFX1 \fadd_0_0_0_0_0/n279_q_reg  ( .D(\fadd_0_0_0_0_0/selectclosepath_d1 ), 
        .CLK(clk), .Q(n13648), .QN(n12838) );
  DFFX1 \fadd_0_0_0_0_2/n279_q_reg  ( .D(\fadd_0_0_0_0_2/selectclosepath_d1 ), 
        .CLK(clk), .Q(n13645), .QN(n12840) );
  DFFX1 \fadd_0_0_0_0_4/n279_q_reg  ( .D(\fadd_0_0_0_0_4/selectclosepath_d1 ), 
        .CLK(clk), .Q(n13644), .QN(n12842) );
  DFFX1 \fadd_0_0_0_0_8/n279_q_reg  ( .D(\fadd_0_0_0_0_8/selectclosepath_d1 ), 
        .CLK(clk), .Q(n13643), .QN(n12846) );
  DFFX1 \fadd_0_0_0_0_10/n279_q_reg  ( .D(\fadd_0_0_0_0_10/n302 ), .CLK(clk), 
        .Q(n13527), .QN(n12068) );
  DFFX1 \current_fsm_reg[43]  ( .D(\U4/Z_43 ), .CLK(clk), .Q(n14185), .QN(
        n12827) );
  DFFX1 \current_fsm_reg[46]  ( .D(\U4/Z_46 ), .CLK(clk), .Q(n14162), .QN(
        n11952) );
  DFFX1 \current_fsm_reg[40]  ( .D(\U4/Z_40 ), .CLK(clk), .Q(n14187), .QN(
        n12828) );
  FADDX1 \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_dualsubclose/sub_1_root_add_300/U2_4  ( 
        .A(\fadd_0_0_0_0_10/U29/Z_3 ), .B(n14975), .CI(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_dualsubclose/sub_1_root_add_300/carry[4] ), .CO(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_dualsubclose/sub_1_root_add_300/carry[5] ), .S(\fadd_0_0_0_0_10/U24/DATA1_4 ) );
  INVX0 U5351 ( .INP(\fadd_0_0_0_0_8/add_859/B[1] ), .ZN(n14872) );
  INVX0 U5352 ( .INP(\fadd_0_0_0_0_9/add_859/B[1] ), .ZN(n14893) );
  INVX0 U5353 ( .INP(n14224), .ZN(n14671) );
  INVX0 U5354 ( .INP(n14228), .ZN(n14777) );
  INVX0 U5355 ( .INP(\fadd_0_0_0_0_6/add_859/B[1] ), .ZN(n14819) );
  INVX0 U5356 ( .INP(n14231), .ZN(n14840) );
  INVX0 U5357 ( .INP(n14229), .ZN(n14798) );
  INVX0 U5358 ( .INP(n14226), .ZN(n14724) );
  INVX0 U5359 ( .INP(n14227), .ZN(n14745) );
  INVX0 U5360 ( .INP(\fadd_0_0_0_0_1/add_859/B[1] ), .ZN(n14692) );
  INVX0 U5361 ( .INP(\fadd_0_0_0_0_10/sub_784/carry[4] ), .ZN(n14176) );
  INVX0 U5362 ( .INP(\fmul_0_0_0_0_10/sub_1_root_add_321/carry[5] ), .ZN(
        n14172) );
  OAI22X1 U5363 ( .IN1(n14979), .IN2(n14968), .IN3(
        \fadd_0_0_0_0_10/U27/DATA1_0 ), .IN4(n14965), .QN(n13467) );
  NAND2X1 U5364 ( .IN1(n9055), .IN2(n14215), .QN(n13516) );
  NAND2X1 U5365 ( .IN1(n9129), .IN2(n14187), .QN(n13634) );
  NOR2X0 U5366 ( .IN1(\fadd_0_0_0_0_8/sub_784/carry [4]), .IN2(
        \fadd_0_0_0_0_8/newx_d1 [8]), .QN(n13654) );
  NOR2X0 U5367 ( .IN1(\fadd_0_0_0_0_9/sub_784/carry [4]), .IN2(
        \fadd_0_0_0_0_9/newx_d1 [8]), .QN(n13655) );
  NOR2X0 U5368 ( .IN1(\fadd_0_0_0_0_0/sub_784/carry [4]), .IN2(
        \fadd_0_0_0_0_0/newx_d1 [8]), .QN(n13656) );
  NOR2X0 U5369 ( .IN1(\fadd_0_0_0_0_4/sub_784/carry [4]), .IN2(
        \fadd_0_0_0_0_4/newx_d1 [8]), .QN(n13657) );
  NOR2X0 U5370 ( .IN1(\fadd_0_0_0_0_6/sub_784/carry [4]), .IN2(
        \fadd_0_0_0_0_6/newx_d1 [8]), .QN(n13658) );
  NOR2X0 U5371 ( .IN1(\fadd_0_0_0_0_7/sub_784/carry [4]), .IN2(
        \fadd_0_0_0_0_7/newx_d1 [8]), .QN(n13659) );
  NOR2X0 U5372 ( .IN1(\fadd_0_0_0_0_5/sub_784/carry [4]), .IN2(
        \fadd_0_0_0_0_5/newx_d1 [8]), .QN(n13660) );
  NOR2X0 U5373 ( .IN1(\fadd_0_0_0_0_2/sub_784/carry [4]), .IN2(
        \fadd_0_0_0_0_2/newx_d1 [8]), .QN(n13661) );
  NOR2X0 U5374 ( .IN1(\fadd_0_0_0_0_3/sub_784/carry [4]), .IN2(
        \fadd_0_0_0_0_3/newx_d1 [8]), .QN(n13662) );
  NOR2X0 U5375 ( .IN1(\fadd_0_0_0_0_1/sub_784/carry [4]), .IN2(
        \fadd_0_0_0_0_1/newx_d1 [8]), .QN(n13663) );
  XOR3X1 U5376 ( .IN1(n14853), .IN2(
        \add_0_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[5] ), .IN3(
        \add_0_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [5]), .Q(\fadd_0_0_0_0_8/fracrcloseymx [5]) );
  XOR3X1 U5377 ( .IN1(n14885), .IN2(
        \add_0_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[5] ), .IN3(
        \add_0_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [5]), .Q(\fadd_0_0_0_0_9/fracrcloseymx [5]) );
  XOR3X1 U5378 ( .IN1(n14663), .IN2(
        \add_0_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[5] ), .IN3(
        \add_0_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [5]), .Q(\fadd_0_0_0_0_0/fracrcloseymx [5]) );
  XOR3X1 U5379 ( .IN1(n14758), .IN2(
        \add_0_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[5] ), .IN3(
        \add_0_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [5]), .Q(\fadd_0_0_0_0_4/fracrcloseymx [5]) );
  XOR3X1 U5380 ( .IN1(n14811), .IN2(
        \add_0_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[5] ), .IN3(
        \add_0_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [5]), .Q(\fadd_0_0_0_0_6/fracrcloseymx [5]) );
  XOR3X1 U5381 ( .IN1(n14832), .IN2(
        \add_0_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[5] ), .IN3(
        \add_0_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [5]), .Q(\fadd_0_0_0_0_7/fracrcloseymx [5]) );
  XOR3X1 U5382 ( .IN1(n14790), .IN2(
        \add_0_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[5] ), .IN3(
        \add_0_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [5]), .Q(\fadd_0_0_0_0_5/fracrcloseymx [5]) );
  XOR3X1 U5383 ( .IN1(n14737), .IN2(
        \add_0_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[5] ), .IN3(
        \add_0_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [5]), .Q(\fadd_0_0_0_0_3/fracrcloseymx [5]) );
  XOR3X1 U5384 ( .IN1(n14705), .IN2(
        \add_0_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[5] ), .IN3(
        \add_0_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [5]), .Q(\fadd_0_0_0_0_2/fracrcloseymx [5]) );
  XOR3X1 U5385 ( .IN1(n14684), .IN2(
        \add_0_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[5] ), .IN3(
        \add_0_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [5]), .Q(\fadd_0_0_0_0_1/fracrcloseymx [5]) );
  NAND2X1 U5386 ( .IN1(n9166), .IN2(n14912), .QN(n14108) );
  INVX0 U5387 ( .INP(rst), .ZN(n14440) );
  NBUFFX2 U5388 ( .INP(n8886), .Z(n14427) );
  NBUFFX2 U5389 ( .INP(n8886), .Z(n14424) );
  NBUFFX2 U5390 ( .INP(n8886), .Z(n14425) );
  NBUFFX2 U5391 ( .INP(n8886), .Z(n14426) );
  NBUFFX2 U5392 ( .INP(n8886), .Z(n14423) );
  NBUFFX2 U5393 ( .INP(n8886), .Z(n14422) );
  INVX0 U5394 ( .INP(n14111), .ZN(n14644) );
  INVX0 U5395 ( .INP(n14110), .ZN(n14647) );
  INVX0 U5396 ( .INP(n14112), .ZN(n14643) );
  INVX0 U5397 ( .INP(n14113), .ZN(n14641) );
  INVX0 U5398 ( .INP(n14109), .ZN(n14648) );
  INVX0 U5399 ( .INP(n14114), .ZN(n14649) );
  INVX0 U5400 ( .INP(n14116), .ZN(n14645) );
  INVX0 U5401 ( .INP(n14115), .ZN(n14646) );
  INVX0 U5402 ( .INP(n14117), .ZN(n14642) );
  NAND2X1 U5403 ( .IN1(n14876), .IN2(n14878), .QN(n10627) );
  NAND2X1 U5404 ( .IN1(n14823), .IN2(n14825), .QN(n10791) );
  NAND2X1 U5405 ( .IN1(n14749), .IN2(n14751), .QN(n11034) );
  NAND2X1 U5406 ( .IN1(n14781), .IN2(n14783), .QN(n10953) );
  NAND2X1 U5407 ( .IN1(n14728), .IN2(n14730), .QN(n11115) );
  NAND2X1 U5408 ( .IN1(n14675), .IN2(n14677), .QN(n11332) );
  NBUFFX2 U5409 ( .INP(n14905), .Z(n14242) );
  NBUFFX2 U5410 ( .INP(n14234), .Z(n14246) );
  NBUFFX2 U5411 ( .INP(n14250), .Z(n14243) );
  NBUFFX2 U5412 ( .INP(n14250), .Z(n14245) );
  NBUFFX2 U5413 ( .INP(n14250), .Z(n14244) );
  NBUFFX2 U5414 ( .INP(n14250), .Z(n14249) );
  NBUFFX2 U5415 ( .INP(n14250), .Z(n14248) );
  NBUFFX2 U5416 ( .INP(n14905), .Z(n14247) );
  NBUFFX2 U5417 ( .INP(n14250), .Z(n14238) );
  NBUFFX2 U5418 ( .INP(n14905), .Z(n14240) );
  NBUFFX2 U5419 ( .INP(n14234), .Z(n14237) );
  NBUFFX2 U5420 ( .INP(n14905), .Z(n14239) );
  NBUFFX2 U5421 ( .INP(n14234), .Z(n14241) );
  NOR2X0 U5422 ( .IN1(n14183), .IN2(n14434), .QN(n8886) );
  NBUFFX2 U5423 ( .INP(n8768), .Z(n14428) );
  NBUFFX2 U5424 ( .INP(n8768), .Z(n14429) );
  NBUFFX2 U5425 ( .INP(n8768), .Z(n14430) );
  NBUFFX2 U5426 ( .INP(n8768), .Z(n14431) );
  NBUFFX2 U5427 ( .INP(n8768), .Z(n14432) );
  INVX0 U5428 ( .INP(n11927), .ZN(n14255) );
  INVX0 U5429 ( .INP(n14435), .ZN(n14433) );
  NAND2X1 U5430 ( .IN1(n14907), .IN2(n14912), .QN(n8674) );
  INVX0 U5431 ( .INP(n14108), .ZN(n14415) );
  INVX0 U5432 ( .INP(n14108), .ZN(n14416) );
  INVX0 U5433 ( .INP(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_dualsubclose/sub_1_root_add_300/carry[5] ), .ZN(n14181) );
  NAND2X1 U5434 ( .IN1(n14939), .IN2(n14963), .QN(n11277) );
  NOR2X0 U5435 ( .IN1(n11442), .IN2(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [5]), .QN(n14109) );
  NOR2X0 U5436 ( .IN1(n11061), .IN2(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [5]), .QN(n14110) );
  NOR2X0 U5437 ( .IN1(n10980), .IN2(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [5]), .QN(n14111) );
  NOR2X0 U5438 ( .IN1(n11223), .IN2(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [5]), .QN(n14112) );
  NOR2X0 U5439 ( .IN1(n11359), .IN2(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [5]), .QN(n14113) );
  INVX0 U5440 ( .INP(n14118), .ZN(n14650) );
  NOR2X0 U5441 ( .IN1(n10654), .IN2(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [5]), .QN(n14114) );
  NOR2X0 U5442 ( .IN1(n10899), .IN2(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [5]), .QN(n14115) );
  NOR2X0 U5443 ( .IN1(n10818), .IN2(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [5]), .QN(n14116) );
  NOR2X0 U5444 ( .IN1(n11142), .IN2(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [5]), .QN(n14117) );
  NOR2X0 U5445 ( .IN1(n10507), .IN2(n14923), .QN(n10502) );
  NOR2X0 U5446 ( .IN1(n14870), .IN2(\fadd_0_0_0_0_8/add_859/B[1] ), .QN(n10673) );
  NOR2X0 U5447 ( .IN1(n14775), .IN2(n14228), .QN(n10999) );
  NOR2X0 U5448 ( .IN1(n14722), .IN2(n14226), .QN(n11161) );
  NOR2X0 U5449 ( .IN1(n14669), .IN2(n14224), .QN(n11378) );
  NOR2X0 U5450 ( .IN1(n14817), .IN2(\fadd_0_0_0_0_6/add_859/B[1] ), .QN(n10837) );
  NOR2X0 U5451 ( .IN1(n14838), .IN2(n14231), .QN(n10756) );
  NOR2X0 U5452 ( .IN1(n14796), .IN2(n14229), .QN(n10918) );
  NOR2X0 U5453 ( .IN1(n14891), .IN2(\fadd_0_0_0_0_9/add_859/B[1] ), .QN(n10592) );
  NOR2X0 U5454 ( .IN1(n14743), .IN2(n14227), .QN(n11080) );
  NOR2X0 U5455 ( .IN1(n14690), .IN2(\fadd_0_0_0_0_1/add_859/B[1] ), .QN(n11297) );
  INVX0 U5456 ( .INP(n12769), .ZN(n14846) );
  NAND2X1 U5457 ( .IN1(n14844), .IN2(n14846), .QN(n10710) );
  INVX0 U5458 ( .INP(n12691), .ZN(n14656) );
  INVX0 U5459 ( .INP(n12751), .ZN(n14804) );
  INVX0 U5460 ( .INP(n12711), .ZN(n14698) );
  INVX0 U5461 ( .INP(n12779), .ZN(n14878) );
  INVX0 U5462 ( .INP(n12731), .ZN(n14751) );
  INVX0 U5463 ( .INP(n12719), .ZN(n14730) );
  INVX0 U5464 ( .INP(n12699), .ZN(n14677) );
  INVX0 U5465 ( .INP(n12759), .ZN(n14825) );
  INVX0 U5466 ( .INP(n12739), .ZN(n14783) );
  NAND2X1 U5467 ( .IN1(n14654), .IN2(n14656), .QN(n11415) );
  NAND2X1 U5468 ( .IN1(n14802), .IN2(n14804), .QN(n10872) );
  NAND2X1 U5469 ( .IN1(n14696), .IN2(n14698), .QN(n11196) );
  INVX0 U5470 ( .INP(n12782), .ZN(n14879) );
  INVX0 U5471 ( .INP(n12762), .ZN(n14826) );
  INVX0 U5472 ( .INP(n12722), .ZN(n14731) );
  INVX0 U5473 ( .INP(n12734), .ZN(n14752) );
  INVX0 U5474 ( .INP(n12742), .ZN(n14784) );
  INVX0 U5475 ( .INP(n12702), .ZN(n14678) );
  INVX0 U5476 ( .INP(n10727), .ZN(n14843) );
  INVX0 U5477 ( .INP(n10644), .ZN(n14875) );
  INVX0 U5478 ( .INP(n10808), .ZN(n14822) );
  INVX0 U5479 ( .INP(n11432), .ZN(n14653) );
  INVX0 U5480 ( .INP(n11051), .ZN(n14748) );
  INVX0 U5481 ( .INP(n10889), .ZN(n14801) );
  INVX0 U5482 ( .INP(n10970), .ZN(n14780) );
  INVX0 U5483 ( .INP(n11132), .ZN(n14727) );
  INVX0 U5484 ( .INP(n11213), .ZN(n14695) );
  INVX0 U5485 ( .INP(n11349), .ZN(n14674) );
  NBUFFX2 U5486 ( .INP(n14905), .Z(n14250) );
  INVX0 U5487 ( .INP(n10715), .ZN(n14844) );
  INVX0 U5488 ( .INP(n11420), .ZN(n14654) );
  INVX0 U5489 ( .INP(n10877), .ZN(n14802) );
  INVX0 U5490 ( .INP(n11201), .ZN(n14696) );
  INVX0 U5491 ( .INP(n10632), .ZN(n14876) );
  INVX0 U5492 ( .INP(n10796), .ZN(n14823) );
  INVX0 U5493 ( .INP(n11039), .ZN(n14749) );
  INVX0 U5494 ( .INP(n10958), .ZN(n14781) );
  INVX0 U5495 ( .INP(n11120), .ZN(n14728) );
  INVX0 U5496 ( .INP(n11337), .ZN(n14675) );
  NBUFFX2 U5497 ( .INP(n14905), .Z(n14236) );
  NBUFFX2 U5498 ( .INP(n14250), .Z(n14235) );
  INVX0 U5499 ( .INP(n11241), .ZN(n14977) );
  INVX0 U5500 ( .INP(n11234), .ZN(n14973) );
  INVX0 U5501 ( .INP(n14279), .ZN(n14276) );
  INVX0 U5502 ( .INP(n14298), .ZN(n14295) );
  INVX0 U5503 ( .INP(n14280), .ZN(n14274) );
  INVX0 U5504 ( .INP(n14299), .ZN(n14293) );
  INVX0 U5505 ( .INP(n14280), .ZN(n14275) );
  INVX0 U5506 ( .INP(n14299), .ZN(n14294) );
  INVX0 U5507 ( .INP(n11927), .ZN(n14254) );
  INVX0 U5508 ( .INP(n8716), .ZN(n14907) );
  INVX0 U5509 ( .INP(n9130), .ZN(n14251) );
  INVX0 U5510 ( .INP(n8679), .ZN(n14909) );
  INVX0 U5511 ( .INP(n8673), .ZN(n14908) );
  INVX0 U5512 ( .INP(n9130), .ZN(n14252) );
  INVX0 U5513 ( .INP(n9130), .ZN(n14253) );
  NBUFFX2 U5514 ( .INP(n14406), .Z(n14413) );
  NBUFFX2 U5515 ( .INP(n14406), .Z(n14412) );
  NBUFFX2 U5516 ( .INP(n9440), .Z(n14411) );
  NBUFFX2 U5517 ( .INP(n14406), .Z(n14409) );
  NBUFFX2 U5518 ( .INP(n9440), .Z(n14408) );
  NBUFFX2 U5519 ( .INP(n9440), .Z(n14407) );
  NBUFFX2 U5520 ( .INP(n14406), .Z(n14410) );
  NOR2X0 U5521 ( .IN1(n14437), .IN2(n14300), .QN(\U4/Z_40 ) );
  NOR2X0 U5522 ( .IN1(n14438), .IN2(n14281), .QN(\U4/Z_36 ) );
  NOR2X0 U5523 ( .IN1(n14438), .IN2(n12829), .QN(\U4/Z_37 ) );
  NOR2X0 U5524 ( .IN1(n14439), .IN2(n11927), .QN(\U4/Z_22 ) );
  INVX0 U5525 ( .INP(n11928), .ZN(n14199) );
  INVX0 U5526 ( .INP(n11928), .ZN(n14198) );
  INVX0 U5527 ( .INP(n11928), .ZN(n14196) );
  INVX0 U5528 ( .INP(n11928), .ZN(n14195) );
  INVX0 U5529 ( .INP(n11928), .ZN(n14194) );
  INVX0 U5530 ( .INP(n11928), .ZN(n14197) );
  INVX0 U5531 ( .INP(n11928), .ZN(n14200) );
  INVX0 U5532 ( .INP(n9410), .ZN(n14912) );
  INVX0 U5533 ( .INP(n13634), .ZN(n14417) );
  INVX0 U5534 ( .INP(n13634), .ZN(n14418) );
  INVX0 U5535 ( .INP(n13516), .ZN(n14420) );
  INVX0 U5536 ( .INP(n13516), .ZN(n14421) );
  NOR2X0 U5537 ( .IN1(n8850), .IN2(n13412), .QN(n8869) );
  NOR2X0 U5538 ( .IN1(n8861), .IN2(n8862), .QN(n8842) );
  NOR2X0 U5539 ( .IN1(n8831), .IN2(n14991), .QN(n8827) );
  INVX0 U5540 ( .INP(n8874), .ZN(n14989) );
  INVX0 U5541 ( .INP(n13412), .ZN(n14993) );
  INVX0 U5542 ( .INP(\fadd_0_0_0_0_10/U25/Z_2 ), .ZN(n14967) );
  INVX0 U5543 ( .INP(\fadd_0_0_0_0_10/U25/Z_3 ), .ZN(n14970) );
  INVX0 U5544 ( .INP(n12794), .ZN(n14975) );
  NOR2X0 U5545 ( .IN1(n11275), .IN2(n11276), .QN(\fadd_0_0_0_0_10/U23/Z_0 ) );
  NOR4X0 U5546 ( .IN1(n11281), .IN2(n11279), .IN3(\fadd_0_0_0_0_10/U24/Z_2 ), 
        .IN4(\fadd_0_0_0_0_10/U24/Z_1 ), .QN(n11275) );
  INVX0 U5547 ( .INP(\fadd_0_0_0_0_0/fracyclose1 [1]), .ZN(n14509) );
  INVX0 U5548 ( .INP(\fadd_0_0_0_0_0/fracrcloseymx [0]), .ZN(n14508) );
  INVX0 U5549 ( .INP(\fadd_0_0_0_0_2/fracyclose1 [1]), .ZN(n14464) );
  INVX0 U5550 ( .INP(\fadd_0_0_0_0_2/fracrcloseymx [0]), .ZN(n14463) );
  INVX0 U5551 ( .INP(\fadd_0_0_0_0_4/fracyclose1 [1]), .ZN(n14500) );
  INVX0 U5552 ( .INP(\fadd_0_0_0_0_4/fracrcloseymx [0]), .ZN(n14499) );
  INVX0 U5553 ( .INP(\fadd_0_0_0_0_5/fracyclose1 [1]), .ZN(n14473) );
  INVX0 U5554 ( .INP(\fadd_0_0_0_0_5/fracrcloseymx [0]), .ZN(n14472) );
  INVX0 U5555 ( .INP(\fadd_0_0_0_0_1/fracyclose1 [1]), .ZN(n14446) );
  INVX0 U5556 ( .INP(\fadd_0_0_0_0_1/fracrcloseymx [0]), .ZN(n14445) );
  INVX0 U5557 ( .INP(\fadd_0_0_0_0_0/fracyclose1 [3]), .ZN(n14512) );
  INVX0 U5558 ( .INP(\fadd_0_0_0_0_0/fracyclose1 [2]), .ZN(n14510) );
  INVX0 U5559 ( .INP(\fadd_0_0_0_0_4/fracyclose1 [3]), .ZN(n14503) );
  INVX0 U5560 ( .INP(\fadd_0_0_0_0_4/fracyclose1 [2]), .ZN(n14501) );
  INVX0 U5561 ( .INP(\fadd_0_0_0_0_5/fracyclose1 [3]), .ZN(n14476) );
  INVX0 U5562 ( .INP(\fadd_0_0_0_0_5/fracyclose1 [2]), .ZN(n14474) );
  INVX0 U5563 ( .INP(\fadd_0_0_0_0_2/fracyclose1 [3]), .ZN(n14467) );
  INVX0 U5564 ( .INP(\fadd_0_0_0_0_2/fracyclose1 [2]), .ZN(n14465) );
  INVX0 U5565 ( .INP(\fadd_0_0_0_0_1/fracyclose1 [3]), .ZN(n14449) );
  INVX0 U5566 ( .INP(\fadd_0_0_0_0_1/fracyclose1 [2]), .ZN(n14447) );
  INVX0 U5567 ( .INP(\fadd_0_0_0_0_0/fracyclose1 [4]), .ZN(n14511) );
  INVX0 U5568 ( .INP(\fadd_0_0_0_0_4/fracyclose1 [4]), .ZN(n14502) );
  INVX0 U5569 ( .INP(\fadd_0_0_0_0_5/fracyclose1 [4]), .ZN(n14475) );
  INVX0 U5570 ( .INP(\fadd_0_0_0_0_2/fracyclose1 [4]), .ZN(n14466) );
  INVX0 U5571 ( .INP(\fadd_0_0_0_0_1/fracyclose1 [4]), .ZN(n14448) );
  NOR2X0 U5572 ( .IN1(n10737), .IN2(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [5]), .QN(n14118) );
  INVX0 U5573 ( .INP(\fadd_0_0_0_0_6/fracyclose1 [1]), .ZN(n14491) );
  INVX0 U5574 ( .INP(\fadd_0_0_0_0_6/fracrcloseymx [0]), .ZN(n14490) );
  INVX0 U5575 ( .INP(\fadd_0_0_0_0_9/fracyclose1 [1]), .ZN(n14518) );
  INVX0 U5576 ( .INP(\fadd_0_0_0_0_9/fracrcloseymx [0]), .ZN(n14517) );
  INVX0 U5577 ( .INP(\fadd_0_0_0_0_7/fracyclose1 [1]), .ZN(n14482) );
  INVX0 U5578 ( .INP(\fadd_0_0_0_0_7/fracrcloseymx [0]), .ZN(n14481) );
  INVX0 U5579 ( .INP(\fadd_0_0_0_0_3/fracyclose1 [1]), .ZN(n14455) );
  INVX0 U5580 ( .INP(\fadd_0_0_0_0_3/fracrcloseymx [0]), .ZN(n14454) );
  INVX0 U5581 ( .INP(\fadd_0_0_0_0_9/fracyclose1 [3]), .ZN(n14521) );
  INVX0 U5582 ( .INP(\fadd_0_0_0_0_6/fracyclose1 [3]), .ZN(n14494) );
  INVX0 U5583 ( .INP(\fadd_0_0_0_0_7/fracyclose1 [3]), .ZN(n14485) );
  INVX0 U5584 ( .INP(\fadd_0_0_0_0_3/fracyclose1 [3]), .ZN(n14458) );
  INVX0 U5585 ( .INP(\fadd_0_0_0_0_9/fracyclose1 [4]), .ZN(n14520) );
  INVX0 U5586 ( .INP(\fadd_0_0_0_0_6/fracyclose1 [4]), .ZN(n14493) );
  INVX0 U5587 ( .INP(\fadd_0_0_0_0_7/fracyclose1 [4]), .ZN(n14484) );
  INVX0 U5588 ( .INP(\fadd_0_0_0_0_3/fracyclose1 [4]), .ZN(n14457) );
  FADDX1 U5589 ( .A(
        \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ), .B(
        n14519), .CI(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [2]), .CO(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [3]), .S(\fadd_0_0_0_0_9/fracrclosexmy [2]) );
  INVX0 U5590 ( .INP(\fadd_0_0_0_0_9/fracyclose1 [2]), .ZN(n14519) );
  FADDX1 U5591 ( .A(
        \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ), .B(
        n14492), .CI(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [2]), .CO(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [3]), .S(\fadd_0_0_0_0_6/fracrclosexmy [2]) );
  INVX0 U5592 ( .INP(\fadd_0_0_0_0_6/fracyclose1 [2]), .ZN(n14492) );
  FADDX1 U5593 ( .A(
        \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ), .B(
        n14483), .CI(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [2]), .CO(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [3]), .S(\fadd_0_0_0_0_7/fracrclosexmy [2]) );
  INVX0 U5594 ( .INP(\fadd_0_0_0_0_7/fracyclose1 [2]), .ZN(n14483) );
  FADDX1 U5595 ( .A(
        \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ), .B(
        n14456), .CI(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [2]), .CO(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [3]), .S(\fadd_0_0_0_0_3/fracrclosexmy [2]) );
  INVX0 U5596 ( .INP(\fadd_0_0_0_0_3/fracyclose1 [2]), .ZN(n14456) );
  OR4X1 U5597 ( .IN1(\fadd_0_0_0_0_8/fracrclosexmy [3]), .IN2(
        \fadd_0_0_0_0_8/fracrclosexmy [4]), .IN3(
        \fadd_0_0_0_0_8/fracrclosexmy [5]), .IN4(n14118), .Q(n10686) );
  OR4X1 U5598 ( .IN1(\fadd_0_0_0_0_9/fracrclosexmy [3]), .IN2(
        \fadd_0_0_0_0_9/fracrclosexmy [4]), .IN3(
        \fadd_0_0_0_0_9/fracrclosexmy [5]), .IN4(n14114), .Q(n10605) );
  OR4X1 U5599 ( .IN1(\fadd_0_0_0_0_6/fracrclosexmy [3]), .IN2(
        \fadd_0_0_0_0_6/fracrclosexmy [4]), .IN3(
        \fadd_0_0_0_0_6/fracrclosexmy [5]), .IN4(n14115), .Q(n10850) );
  OR4X1 U5600 ( .IN1(\fadd_0_0_0_0_7/fracrclosexmy [3]), .IN2(
        \fadd_0_0_0_0_7/fracrclosexmy [4]), .IN3(
        \fadd_0_0_0_0_7/fracrclosexmy [5]), .IN4(n14116), .Q(n10769) );
  OR4X1 U5601 ( .IN1(\fadd_0_0_0_0_3/fracrclosexmy [3]), .IN2(
        \fadd_0_0_0_0_3/fracrclosexmy [4]), .IN3(
        \fadd_0_0_0_0_3/fracrclosexmy [5]), .IN4(n14117), .Q(n11093) );
  INVX0 U5602 ( .INP(n8826), .ZN(n14988) );
  OR4X1 U5603 ( .IN1(\fadd_0_0_0_0_0/fracrclosexmy [3]), .IN2(
        \fadd_0_0_0_0_0/fracrclosexmy [4]), .IN3(
        \fadd_0_0_0_0_0/fracrclosexmy [5]), .IN4(n14109), .Q(n11391) );
  OR4X1 U5604 ( .IN1(\fadd_0_0_0_0_4/fracrclosexmy [3]), .IN2(
        \fadd_0_0_0_0_4/fracrclosexmy [4]), .IN3(
        \fadd_0_0_0_0_4/fracrclosexmy [5]), .IN4(n14110), .Q(n11012) );
  OR4X1 U5605 ( .IN1(\fadd_0_0_0_0_5/fracrclosexmy [3]), .IN2(
        \fadd_0_0_0_0_5/fracrclosexmy [4]), .IN3(
        \fadd_0_0_0_0_5/fracrclosexmy [5]), .IN4(n14111), .Q(n10931) );
  OR4X1 U5606 ( .IN1(\fadd_0_0_0_0_2/fracrclosexmy [3]), .IN2(
        \fadd_0_0_0_0_2/fracrclosexmy [4]), .IN3(
        \fadd_0_0_0_0_2/fracrclosexmy [5]), .IN4(n14112), .Q(n11174) );
  OR4X1 U5607 ( .IN1(\fadd_0_0_0_0_1/fracrclosexmy [3]), .IN2(
        \fadd_0_0_0_0_1/fracrclosexmy [4]), .IN3(
        \fadd_0_0_0_0_1/fracrclosexmy [5]), .IN4(n14113), .Q(n11310) );
  OR3X1 U5608 ( .IN1(\fadd_0_0_0_0_0/fracrcloseymx [0]), .IN2(
        \fadd_0_0_0_0_0/fracrcloseymx [1]), .IN3(n11396), .Q(n11394) );
  OR3X1 U5609 ( .IN1(\fadd_0_0_0_0_4/fracrcloseymx [0]), .IN2(
        \fadd_0_0_0_0_4/fracrcloseymx [1]), .IN3(n11017), .Q(n11015) );
  OR3X1 U5610 ( .IN1(\fadd_0_0_0_0_5/fracrcloseymx [0]), .IN2(
        \fadd_0_0_0_0_5/fracrcloseymx [1]), .IN3(n10936), .Q(n10934) );
  OR3X1 U5611 ( .IN1(\fadd_0_0_0_0_2/fracrcloseymx [0]), .IN2(
        \fadd_0_0_0_0_2/fracrcloseymx [1]), .IN3(n11179), .Q(n11177) );
  OR3X1 U5612 ( .IN1(\fadd_0_0_0_0_1/fracrcloseymx [0]), .IN2(
        \fadd_0_0_0_0_1/fracrcloseymx [1]), .IN3(n11315), .Q(n11313) );
  INVX0 U5613 ( .INP(n10487), .ZN(n14920) );
  NAND2X1 U5614 ( .IN1(n14174), .IN2(n14175), .QN(
        \fmul_0_0_0_0_10/sub_1_root_add_321/carry[5] ) );
  INVX0 U5615 ( .INP(n14122), .ZN(n14174) );
  AND2X1 U5616 ( .IN1(n14172), .IN2(n14173), .Q(n14119) );
  NAND2X1 U5617 ( .IN1(n10549), .IN2(n10548), .QN(n10494) );
  INVX0 U5618 ( .INP(n10548), .ZN(n14927) );
  INVX0 U5619 ( .INP(n10549), .ZN(n14926) );
  INVX0 U5620 ( .INP(\fadd_0_0_0_0_10/U29/Z_1 ), .ZN(n14966) );
  NAND2X1 U5621 ( .IN1(\fadd_0_0_0_0_10/U29/Z_0 ), .IN2(n13467), .QN(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_dualsubclose/sub_1_root_add_303/carry[2] ) );
  INVX0 U5622 ( .INP(\fadd_0_0_0_0_10/U29/Z_2 ), .ZN(n14969) );
  INVX0 U5623 ( .INP(\fadd_0_0_0_0_10/U29/Z_3 ), .ZN(n14972) );
  INVX0 U5624 ( .INP(
        \add_0_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .ZN(n14504) );
  INVX0 U5625 ( .INP(
        \add_0_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .ZN(n14486) );
  INVX0 U5626 ( .INP(
        \add_0_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .ZN(n14459) );
  INVX0 U5627 ( .INP(
        \add_0_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .ZN(n14513) );
  INVX0 U5628 ( .INP(
        \add_0_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .ZN(n14495) );
  INVX0 U5629 ( .INP(
        \add_0_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .ZN(n14477) );
  INVX0 U5630 ( .INP(
        \add_0_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .ZN(n14468) );
  INVX0 U5631 ( .INP(
        \add_0_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .ZN(n14450) );
  INVX0 U5632 ( .INP(
        \add_0_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .ZN(n14441) );
  NBUFFX2 U5633 ( .INP(\fadd_0_0_0_0_4/add_859/B[1] ), .Z(n14228) );
  NBUFFX2 U5634 ( .INP(\fadd_0_0_0_0_2/add_859/B[1] ), .Z(n14226) );
  INVX0 U5635 ( .INP(\fadd_0_0_0_0_10/U29/Z_0 ), .ZN(n14962) );
  INVX0 U5636 ( .INP(
        \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ), .ZN(
        n14487) );
  INVX0 U5637 ( .INP(
        \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ), .ZN(
        n14514) );
  INVX0 U5638 ( .INP(
        \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ), .ZN(
        n14478) );
  INVX0 U5639 ( .INP(
        \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ), .ZN(
        n14451) );
  INVX0 U5640 ( .INP(
        \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ), .ZN(
        n14505) );
  INVX0 U5641 ( .INP(
        \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ), .ZN(
        n14460) );
  INVX0 U5642 ( .INP(
        \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ), .ZN(
        n14496) );
  INVX0 U5643 ( .INP(
        \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ), .ZN(
        n14469) );
  INVX0 U5644 ( .INP(
        \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ), .ZN(
        n14442) );
  INVX0 U5645 ( .INP(n10539), .ZN(n14925) );
  NBUFFX2 U5646 ( .INP(\fadd_0_0_0_0_8/add_859/B[1] ), .Z(n14232) );
  INVX0 U5647 ( .INP(n10510), .ZN(n14923) );
  INVX0 U5648 ( .INP(
        \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ), .ZN(
        n14506) );
  INVX0 U5649 ( .INP(
        \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ), .ZN(
        n14488) );
  INVX0 U5650 ( .INP(
        \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ), .ZN(
        n14461) );
  INVX0 U5651 ( .INP(
        \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ), .ZN(
        n14515) );
  INVX0 U5652 ( .INP(
        \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ), .ZN(
        n14497) );
  INVX0 U5653 ( .INP(
        \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ), .ZN(
        n14479) );
  INVX0 U5654 ( .INP(
        \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ), .ZN(
        n14470) );
  INVX0 U5655 ( .INP(
        \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ), .ZN(
        n14452) );
  INVX0 U5656 ( .INP(
        \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ), .ZN(
        n14443) );
  NBUFFX2 U5657 ( .INP(\fadd_0_0_0_0_0/add_859/B[1] ), .Z(n14224) );
  NBUFFX2 U5658 ( .INP(\fadd_0_0_0_0_7/add_859/B[1] ), .Z(n14231) );
  NBUFFX2 U5659 ( .INP(\fadd_0_0_0_0_5/add_859/B[1] ), .Z(n14229) );
  NBUFFX2 U5660 ( .INP(\fadd_0_0_0_0_3/add_859/B[1] ), .Z(n14227) );
  NBUFFX2 U5661 ( .INP(\fadd_0_0_0_0_6/add_859/B[1] ), .Z(n14230) );
  NBUFFX2 U5662 ( .INP(\fadd_0_0_0_0_9/add_859/B[1] ), .Z(n14233) );
  NBUFFX2 U5663 ( .INP(\fadd_0_0_0_0_1/add_859/B[1] ), .Z(n14225) );
  INVX0 U5664 ( .INP(
        \fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ), .ZN(
        n14507) );
  INVX0 U5665 ( .INP(
        \fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ), .ZN(
        n14489) );
  INVX0 U5666 ( .INP(
        \fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ), .ZN(
        n14462) );
  INVX0 U5667 ( .INP(
        \fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ), .ZN(
        n14516) );
  INVX0 U5668 ( .INP(
        \fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ), .ZN(
        n14498) );
  INVX0 U5669 ( .INP(
        \fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ), .ZN(
        n14480) );
  INVX0 U5670 ( .INP(
        \fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ), .ZN(
        n14471) );
  INVX0 U5671 ( .INP(
        \fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ), .ZN(
        n14453) );
  INVX0 U5672 ( .INP(
        \fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ), .ZN(
        n14444) );
  NAND2X1 U5673 ( .IN1(n14853), .IN2(n10735), .QN(n12769) );
  NAND2X1 U5674 ( .IN1(n14663), .IN2(n11440), .QN(n12691) );
  NAND2X1 U5675 ( .IN1(n14811), .IN2(n10897), .QN(n12751) );
  NAND2X1 U5676 ( .IN1(n14705), .IN2(n11221), .QN(n12711) );
  NAND2X1 U5677 ( .IN1(n14885), .IN2(n10652), .QN(n12779) );
  NAND2X1 U5678 ( .IN1(n14758), .IN2(n11059), .QN(n12731) );
  NAND2X1 U5679 ( .IN1(n14832), .IN2(n10816), .QN(n12759) );
  NAND2X1 U5680 ( .IN1(n14790), .IN2(n10978), .QN(n12739) );
  NAND2X1 U5681 ( .IN1(n14737), .IN2(n11140), .QN(n12719) );
  NAND2X1 U5682 ( .IN1(n14684), .IN2(n11357), .QN(n12699) );
  INVX0 U5683 ( .INP(\fadd_0_0_0_0_8/expoperationsel[0] ), .ZN(n14870) );
  INVX0 U5684 ( .INP(\fadd_0_0_0_0_4/expoperationsel[0] ), .ZN(n14775) );
  INVX0 U5685 ( .INP(\fadd_0_0_0_0_2/expoperationsel[0] ), .ZN(n14722) );
  INVX0 U5686 ( .INP(n12772), .ZN(n14847) );
  INVX0 U5687 ( .INP(n10693), .ZN(n14841) );
  INVX0 U5688 ( .INP(n12754), .ZN(n14805) );
  INVX0 U5689 ( .INP(n10612), .ZN(n14873) );
  INVX0 U5690 ( .INP(n10857), .ZN(n14799) );
  INVX0 U5691 ( .INP(n10776), .ZN(n14820) );
  INVX0 U5692 ( .INP(n11100), .ZN(n14725) );
  INVX0 U5693 ( .INP(n12694), .ZN(n14657) );
  INVX0 U5694 ( .INP(n12714), .ZN(n14699) );
  INVX0 U5695 ( .INP(n11398), .ZN(n14651) );
  INVX0 U5696 ( .INP(n11019), .ZN(n14746) );
  INVX0 U5697 ( .INP(n10938), .ZN(n14778) );
  INVX0 U5698 ( .INP(n11181), .ZN(n14693) );
  INVX0 U5699 ( .INP(n11317), .ZN(n14672) );
  NAND2X1 U5700 ( .IN1(n14845), .IN2(n10723), .QN(n10727) );
  INVX0 U5701 ( .INP(n10729), .ZN(n14845) );
  NAND2X1 U5702 ( .IN1(n14655), .IN2(n11428), .QN(n11432) );
  NAND2X1 U5703 ( .IN1(n14803), .IN2(n10885), .QN(n10889) );
  NAND2X1 U5704 ( .IN1(n14697), .IN2(n11209), .QN(n11213) );
  INVX0 U5705 ( .INP(n11434), .ZN(n14655) );
  INVX0 U5706 ( .INP(n10891), .ZN(n14803) );
  INVX0 U5707 ( .INP(n11215), .ZN(n14697) );
  NAND2X1 U5708 ( .IN1(n14877), .IN2(n10640), .QN(n10644) );
  NAND2X1 U5709 ( .IN1(n14824), .IN2(n10804), .QN(n10808) );
  NAND2X1 U5710 ( .IN1(n14750), .IN2(n11047), .QN(n11051) );
  NAND2X1 U5711 ( .IN1(n14782), .IN2(n10966), .QN(n10970) );
  NAND2X1 U5712 ( .IN1(n14729), .IN2(n11128), .QN(n11132) );
  NAND2X1 U5713 ( .IN1(n14676), .IN2(n11345), .QN(n11349) );
  INVX0 U5714 ( .INP(n10646), .ZN(n14877) );
  INVX0 U5715 ( .INP(n11053), .ZN(n14750) );
  INVX0 U5716 ( .INP(n10810), .ZN(n14824) );
  INVX0 U5717 ( .INP(n10972), .ZN(n14782) );
  INVX0 U5718 ( .INP(n11134), .ZN(n14729) );
  INVX0 U5719 ( .INP(n11351), .ZN(n14676) );
  NAND2X1 U5720 ( .IN1(n10729), .IN2(n10723), .QN(n10715) );
  NAND2X1 U5721 ( .IN1(n11434), .IN2(n11428), .QN(n11420) );
  NAND2X1 U5722 ( .IN1(n10891), .IN2(n10885), .QN(n10877) );
  NAND2X1 U5723 ( .IN1(n11215), .IN2(n11209), .QN(n11201) );
  NAND2X1 U5724 ( .IN1(n10646), .IN2(n10640), .QN(n10632) );
  NAND2X1 U5725 ( .IN1(n10810), .IN2(n10804), .QN(n10796) );
  NAND2X1 U5726 ( .IN1(n11053), .IN2(n11047), .QN(n11039) );
  NAND2X1 U5727 ( .IN1(n10972), .IN2(n10966), .QN(n10958) );
  NAND2X1 U5728 ( .IN1(n11134), .IN2(n11128), .QN(n11120) );
  NAND2X1 U5729 ( .IN1(n11351), .IN2(n11345), .QN(n11337) );
  INVX0 U5730 ( .INP(n10723), .ZN(n14842) );
  INVX0 U5731 ( .INP(n11428), .ZN(n14652) );
  INVX0 U5732 ( .INP(n10885), .ZN(n14800) );
  INVX0 U5733 ( .INP(n11209), .ZN(n14694) );
  INVX0 U5734 ( .INP(n10640), .ZN(n14874) );
  INVX0 U5735 ( .INP(n11047), .ZN(n14747) );
  INVX0 U5736 ( .INP(n10804), .ZN(n14821) );
  INVX0 U5737 ( .INP(n10966), .ZN(n14779) );
  INVX0 U5738 ( .INP(n11128), .ZN(n14726) );
  INVX0 U5739 ( .INP(n11345), .ZN(n14673) );
  INVX0 U5740 ( .INP(\fadd_0_0_0_0_0/expoperationsel[0] ), .ZN(n14669) );
  INVX0 U5741 ( .INP(\fadd_0_0_0_0_6/expoperationsel[0] ), .ZN(n14817) );
  INVX0 U5742 ( .INP(\fadd_0_0_0_0_7/expoperationsel[0] ), .ZN(n14838) );
  INVX0 U5743 ( .INP(\fadd_0_0_0_0_5/expoperationsel[0] ), .ZN(n14796) );
  INVX0 U5744 ( .INP(\fadd_0_0_0_0_9/expoperationsel[0] ), .ZN(n14891) );
  INVX0 U5745 ( .INP(\fadd_0_0_0_0_3/expoperationsel[0] ), .ZN(n14743) );
  INVX0 U5746 ( .INP(\fadd_0_0_0_0_1/expoperationsel[0] ), .ZN(n14690) );
  NBUFFX2 U5747 ( .INP(n14905), .Z(n14234) );
  INVX0 U5748 ( .INP(n11279), .ZN(n14939) );
  INVX0 U5749 ( .INP(n13401), .ZN(n14964) );
  INVX0 U5750 ( .INP(n9009), .ZN(n14911) );
  INVX0 U5751 ( .INP(n11242), .ZN(n14978) );
  NBUFFX2 U5752 ( .INP(n14396), .Z(n14405) );
  NBUFFX2 U5753 ( .INP(n14396), .Z(n14404) );
  NBUFFX2 U5754 ( .INP(n14396), .Z(n14403) );
  NBUFFX2 U5755 ( .INP(n14395), .Z(n14402) );
  NBUFFX2 U5756 ( .INP(n14395), .Z(n14401) );
  NBUFFX2 U5757 ( .INP(n14395), .Z(n14400) );
  NBUFFX2 U5758 ( .INP(n9441), .Z(n14399) );
  NBUFFX2 U5759 ( .INP(n14396), .Z(n14398) );
  NBUFFX2 U5760 ( .INP(n14395), .Z(n14397) );
  NAND2X1 U5761 ( .IN1(\fadd_0_0_0_0_10/U27/Z_1 ), .IN2(n14976), .QN(n11252)
         );
  INVX0 U5762 ( .INP(n11240), .ZN(n14938) );
  NBUFFX2 U5763 ( .INP(n14363), .Z(n14355) );
  NBUFFX2 U5764 ( .INP(n14363), .Z(n14356) );
  NBUFFX2 U5765 ( .INP(n14362), .Z(n14357) );
  NBUFFX2 U5766 ( .INP(n14361), .Z(n14358) );
  NBUFFX2 U5767 ( .INP(n14361), .Z(n14359) );
  NBUFFX2 U5768 ( .INP(n9451), .Z(n14345) );
  NBUFFX2 U5769 ( .INP(n9451), .Z(n14346) );
  NBUFFX2 U5770 ( .INP(n14344), .Z(n14347) );
  NBUFFX2 U5771 ( .INP(n14344), .Z(n14348) );
  NBUFFX2 U5772 ( .INP(n14344), .Z(n14349) );
  NBUFFX2 U5773 ( .INP(n14344), .Z(n14350) );
  NBUFFX2 U5774 ( .INP(n14344), .Z(n14351) );
  NBUFFX2 U5775 ( .INP(n14344), .Z(n14352) );
  NBUFFX2 U5776 ( .INP(n14344), .Z(n14353) );
  NBUFFX2 U5777 ( .INP(n14344), .Z(n14354) );
  NBUFFX2 U5778 ( .INP(n14361), .Z(n14360) );
  NBUFFX2 U5779 ( .INP(n9446), .Z(n14376) );
  NBUFFX2 U5780 ( .INP(n9446), .Z(n14377) );
  NBUFFX2 U5781 ( .INP(n14375), .Z(n14378) );
  NBUFFX2 U5782 ( .INP(n14375), .Z(n14379) );
  NBUFFX2 U5783 ( .INP(n14375), .Z(n14380) );
  NBUFFX2 U5784 ( .INP(n14375), .Z(n14381) );
  NBUFFX2 U5785 ( .INP(n14375), .Z(n14382) );
  NBUFFX2 U5786 ( .INP(n14375), .Z(n14383) );
  NBUFFX2 U5787 ( .INP(n14375), .Z(n14384) );
  NBUFFX2 U5788 ( .INP(n14375), .Z(n14385) );
  NBUFFX2 U5789 ( .INP(n9447), .Z(n14364) );
  NBUFFX2 U5790 ( .INP(n9447), .Z(n14365) );
  NBUFFX2 U5791 ( .INP(n14374), .Z(n14366) );
  NBUFFX2 U5792 ( .INP(n9447), .Z(n14367) );
  NBUFFX2 U5793 ( .INP(n14374), .Z(n14368) );
  NBUFFX2 U5794 ( .INP(n9447), .Z(n14369) );
  NBUFFX2 U5795 ( .INP(n9447), .Z(n14370) );
  NBUFFX2 U5796 ( .INP(n14374), .Z(n14371) );
  NBUFFX2 U5797 ( .INP(n14374), .Z(n14372) );
  NBUFFX2 U5798 ( .INP(n14374), .Z(n14373) );
  INVX0 U5799 ( .INP(\fadd_0_0_0_0_9/sub_784/B[1] ), .ZN(n14937) );
  INVX0 U5800 ( .INP(\fadd_0_0_0_0_8/sub_784/B[1] ), .ZN(n14936) );
  INVX0 U5801 ( .INP(\fadd_0_0_0_0_7/sub_784/B[1] ), .ZN(n14935) );
  INVX0 U5802 ( .INP(\fadd_0_0_0_0_6/sub_784/B[1] ), .ZN(n14934) );
  INVX0 U5803 ( .INP(\fadd_0_0_0_0_5/sub_784/B[1] ), .ZN(n14933) );
  INVX0 U5804 ( .INP(\fadd_0_0_0_0_4/sub_784/B[1] ), .ZN(n14932) );
  INVX0 U5805 ( .INP(\fadd_0_0_0_0_3/sub_784/B[1] ), .ZN(n14931) );
  INVX0 U5806 ( .INP(\fadd_0_0_0_0_2/sub_784/B[1] ), .ZN(n14930) );
  INVX0 U5807 ( .INP(\fadd_0_0_0_0_1/sub_784/B[1] ), .ZN(n14929) );
  INVX0 U5808 ( .INP(\fadd_0_0_0_0_0/sub_784/B[1] ), .ZN(n14928) );
  NBUFFX2 U5809 ( .INP(n9452), .Z(n14334) );
  NBUFFX2 U5810 ( .INP(n9452), .Z(n14335) );
  NBUFFX2 U5811 ( .INP(n9452), .Z(n14336) );
  NBUFFX2 U5812 ( .INP(n9452), .Z(n14337) );
  NBUFFX2 U5813 ( .INP(n9452), .Z(n14338) );
  NBUFFX2 U5814 ( .INP(n9452), .Z(n14339) );
  NBUFFX2 U5815 ( .INP(n9452), .Z(n14340) );
  NBUFFX2 U5816 ( .INP(n9452), .Z(n14341) );
  NBUFFX2 U5817 ( .INP(n9452), .Z(n14342) );
  NBUFFX2 U5818 ( .INP(n9452), .Z(n14343) );
  NBUFFX2 U5819 ( .INP(n9454), .Z(n14325) );
  NBUFFX2 U5820 ( .INP(n9454), .Z(n14326) );
  NBUFFX2 U5821 ( .INP(n9454), .Z(n14327) );
  NBUFFX2 U5822 ( .INP(n14324), .Z(n14328) );
  NBUFFX2 U5823 ( .INP(n9454), .Z(n14329) );
  NBUFFX2 U5824 ( .INP(n9454), .Z(n14330) );
  NBUFFX2 U5825 ( .INP(n14324), .Z(n14331) );
  NBUFFX2 U5826 ( .INP(n14324), .Z(n14332) );
  NBUFFX2 U5827 ( .INP(n14324), .Z(n14333) );
  NBUFFX2 U5828 ( .INP(n14323), .Z(n14313) );
  NBUFFX2 U5829 ( .INP(n9455), .Z(n14314) );
  NBUFFX2 U5830 ( .INP(n14323), .Z(n14315) );
  NBUFFX2 U5831 ( .INP(n14323), .Z(n14316) );
  NBUFFX2 U5832 ( .INP(n14323), .Z(n14317) );
  NBUFFX2 U5833 ( .INP(n9455), .Z(n14318) );
  NBUFFX2 U5834 ( .INP(n9455), .Z(n14319) );
  NBUFFX2 U5835 ( .INP(n9455), .Z(n14320) );
  NBUFFX2 U5836 ( .INP(n14323), .Z(n14321) );
  NBUFFX2 U5837 ( .INP(n14323), .Z(n14322) );
  NBUFFX2 U5838 ( .INP(n9443), .Z(n14394) );
  NBUFFX2 U5839 ( .INP(n9443), .Z(n14393) );
  NBUFFX2 U5840 ( .INP(n9443), .Z(n14392) );
  NBUFFX2 U5841 ( .INP(n9443), .Z(n14391) );
  NBUFFX2 U5842 ( .INP(n9443), .Z(n14390) );
  NBUFFX2 U5843 ( .INP(n9443), .Z(n14389) );
  NBUFFX2 U5844 ( .INP(n9443), .Z(n14388) );
  NBUFFX2 U5845 ( .INP(n9443), .Z(n14387) );
  NBUFFX2 U5846 ( .INP(n9443), .Z(n14386) );
  NAND2X1 U5847 ( .IN1(n10422), .IN2(n10423), .QN(\fmul_0_0_0_0_9/round ) );
  NAND2X1 U5848 ( .IN1(n10430), .IN2(n10431), .QN(\fmul_0_0_0_0_8/round ) );
  NAND2X1 U5849 ( .IN1(n10438), .IN2(n10439), .QN(\fmul_0_0_0_0_7/round ) );
  NAND2X1 U5850 ( .IN1(n10446), .IN2(n10447), .QN(\fmul_0_0_0_0_6/round ) );
  NAND2X1 U5851 ( .IN1(n10454), .IN2(n10455), .QN(\fmul_0_0_0_0_5/round ) );
  NAND2X1 U5852 ( .IN1(n10462), .IN2(n10463), .QN(\fmul_0_0_0_0_4/round ) );
  NAND2X1 U5853 ( .IN1(n10470), .IN2(n10471), .QN(\fmul_0_0_0_0_3/round ) );
  NAND2X1 U5854 ( .IN1(n10478), .IN2(n10479), .QN(\fmul_0_0_0_0_2/round ) );
  NAND2X1 U5855 ( .IN1(n10568), .IN2(n10569), .QN(\fmul_0_0_0_0_1/round ) );
  NAND2X1 U5856 ( .IN1(n8764), .IN2(n8763), .QN(n8716) );
  NAND2X1 U5857 ( .IN1(n14215), .IN2(n8763), .QN(n8679) );
  NAND2X0 U5858 ( .IN1(n8763), .IN2(n14187), .QN(n8673) );
  INVX0 U5859 ( .INP(n8680), .ZN(n14906) );
  AO21X1 U5860 ( .IN1(n14240), .IN2(n13498), .IN3(n9436), .Q(n13136) );
  INVX0 U5861 ( .INP(n14440), .ZN(n14437) );
  NOR2X0 U5862 ( .IN1(n14437), .IN2(n13715), .QN(n13442) );
  NOR2X0 U5863 ( .IN1(rst), .IN2(n13476), .QN(\U4/Z_9 ) );
  NOR2X0 U5864 ( .IN1(rst), .IN2(n13631), .QN(n13437) );
  NBUFFX2 U5865 ( .INP(n14406), .Z(n14414) );
  NBUFFX2 U5866 ( .INP(n9440), .Z(n14406) );
  INVX0 U5867 ( .INP(n14137), .ZN(n14215) );
  INVX0 U5868 ( .INP(n14440), .ZN(n14438) );
  INVX0 U5869 ( .INP(n14440), .ZN(n14439) );
  NOR2X0 U5870 ( .IN1(\fadd_0_0_0_0_10/U21/DATA2_3 ), .IN2(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/SUM[7] ), .QN(n13412) );
  NOR2X0 U5871 ( .IN1(n8809), .IN2(n8810), .QN(n8791) );
  NAND2X1 U5872 ( .IN1(n8870), .IN2(n8871), .QN(n8861) );
  NAND2X1 U5873 ( .IN1(n8827), .IN2(n8828), .QN(n8809) );
  INVX0 U5874 ( .INP(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/carry[6] ), .ZN(n14171) );
  NOR2X0 U5875 ( .IN1(n14995), .IN2(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/SUM[7] ), .QN(n8850) );
  INVX0 U5876 ( .INP(\fadd_0_0_0_0_10/U21/DATA2_3 ), .ZN(n14995) );
  INVX0 U5877 ( .INP(n8838), .ZN(n14990) );
  INVX0 U5878 ( .INP(n8805), .ZN(n14994) );
  INVX0 U5879 ( .INP(\fadd_0_0_0_0_10/U27/DATA1_0 ), .ZN(n14979) );
  NAND2X1 U5880 ( .IN1(n14979), .IN2(n14181), .QN(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_dualsubclose/sub_1_root_add_300/carry[6] ) );
  INVX0 U5881 ( .INP(n11255), .ZN(n14968) );
  INVX0 U5882 ( .INP(n11262), .ZN(n14965) );
  NAND2X1 U5883 ( .IN1(\fadd_0_0_0_0_10/U27/DATA1_0 ), .IN2(n14965), .QN(
        n13401) );
  INVX0 U5884 ( .INP(n11442), .ZN(n14663) );
  INVX0 U5885 ( .INP(n11223), .ZN(n14705) );
  INVX0 U5886 ( .INP(n11061), .ZN(n14758) );
  INVX0 U5887 ( .INP(n10980), .ZN(n14790) );
  INVX0 U5888 ( .INP(n11359), .ZN(n14684) );
  NOR2X0 U5889 ( .IN1(n14663), .IN2(n11443), .QN(
        \fadd_0_0_0_0_0/fracrcloseymx [0]) );
  NOR2X0 U5890 ( .IN1(n14758), .IN2(n11062), .QN(
        \fadd_0_0_0_0_4/fracrcloseymx [0]) );
  NOR2X0 U5891 ( .IN1(n14790), .IN2(n10981), .QN(
        \fadd_0_0_0_0_5/fracrcloseymx [0]) );
  NOR2X0 U5892 ( .IN1(n14705), .IN2(n11224), .QN(
        \fadd_0_0_0_0_2/fracrcloseymx [0]) );
  NOR2X0 U5893 ( .IN1(n14684), .IN2(n11360), .QN(
        \fadd_0_0_0_0_1/fracrcloseymx [0]) );
  INVX0 U5894 ( .INP(n10737), .ZN(n14853) );
  NOR2X0 U5895 ( .IN1(n14853), .IN2(n10738), .QN(
        \fadd_0_0_0_0_8/fracrcloseymx [0]) );
  INVX0 U5896 ( .INP(\fadd_0_0_0_0_8/fracyclose1 [1]), .ZN(n14527) );
  INVX0 U5897 ( .INP(\fadd_0_0_0_0_8/fracrcloseymx [0]), .ZN(n14526) );
  INVX0 U5898 ( .INP(\fadd_0_0_0_0_8/fracyclose1 [3]), .ZN(n14530) );
  INVX0 U5899 ( .INP(\fadd_0_0_0_0_8/fracyclose1 [4]), .ZN(n14529) );
  FADDX1 U5900 ( .A(
        \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ), .B(
        n14528), .CI(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [2]), .CO(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [3]), .S(\fadd_0_0_0_0_8/fracrclosexmy [2]) );
  INVX0 U5901 ( .INP(\fadd_0_0_0_0_8/fracyclose1 [2]), .ZN(n14528) );
  INVX0 U5902 ( .INP(n10899), .ZN(n14811) );
  INVX0 U5903 ( .INP(n10654), .ZN(n14885) );
  INVX0 U5904 ( .INP(n10818), .ZN(n14832) );
  INVX0 U5905 ( .INP(n11142), .ZN(n14737) );
  NOR2X0 U5906 ( .IN1(n14885), .IN2(n10655), .QN(
        \fadd_0_0_0_0_9/fracrcloseymx [0]) );
  NOR2X0 U5907 ( .IN1(n14811), .IN2(n10900), .QN(
        \fadd_0_0_0_0_6/fracrcloseymx [0]) );
  NOR2X0 U5908 ( .IN1(n14832), .IN2(n10819), .QN(
        \fadd_0_0_0_0_7/fracrcloseymx [0]) );
  NOR2X0 U5909 ( .IN1(n14737), .IN2(n11143), .QN(
        \fadd_0_0_0_0_3/fracrcloseymx [0]) );
  NOR2X0 U5910 ( .IN1(n13677), .IN2(n8839), .QN(n11268) );
  XOR2X1 U5911 ( .IN1(n11396), .IN2(n11397), .Q(n11395) );
  XOR2X1 U5912 ( .IN1(n11017), .IN2(n11018), .Q(n11016) );
  XOR2X1 U5913 ( .IN1(n10936), .IN2(n10937), .Q(n10935) );
  XOR2X1 U5914 ( .IN1(n11179), .IN2(n11180), .Q(n11178) );
  XOR2X1 U5915 ( .IN1(n11315), .IN2(n11316), .Q(n11314) );
  INVX0 U5916 ( .INP(n8804), .ZN(n14987) );
  NAND2X1 U5917 ( .IN1(n8839), .IN2(n13677), .QN(n8837) );
  INVX0 U5918 ( .INP(n11443), .ZN(n14662) );
  INVX0 U5919 ( .INP(n11224), .ZN(n14704) );
  INVX0 U5920 ( .INP(n11062), .ZN(n14757) );
  INVX0 U5921 ( .INP(n10981), .ZN(n14789) );
  INVX0 U5922 ( .INP(n11360), .ZN(n14683) );
  INVX0 U5923 ( .INP(n10738), .ZN(n14852) );
  INVX0 U5924 ( .INP(n10900), .ZN(n14810) );
  INVX0 U5925 ( .INP(n10655), .ZN(n14884) );
  INVX0 U5926 ( .INP(n10819), .ZN(n14831) );
  INVX0 U5927 ( .INP(n11143), .ZN(n14736) );
  INVX0 U5928 ( .INP(n11433), .ZN(n14661) );
  INVX0 U5929 ( .INP(n11214), .ZN(n14703) );
  INVX0 U5930 ( .INP(n11052), .ZN(n14756) );
  INVX0 U5931 ( .INP(n10971), .ZN(n14788) );
  INVX0 U5932 ( .INP(n11350), .ZN(n14682) );
  INVX0 U5933 ( .INP(n10728), .ZN(n14851) );
  INVX0 U5934 ( .INP(n10890), .ZN(n14809) );
  INVX0 U5935 ( .INP(n10645), .ZN(n14883) );
  INVX0 U5936 ( .INP(n10809), .ZN(n14830) );
  INVX0 U5937 ( .INP(n11133), .ZN(n14735) );
  INVX0 U5938 ( .INP(n11251), .ZN(n14971) );
  INVX0 U5939 ( .INP(n8844), .ZN(n14991) );
  NOR2X0 U5940 ( .IN1(n10562), .IN2(n10563), .QN(n10561) );
  NAND2X1 U5941 ( .IN1(n13618), .IN2(n13468), .QN(n10558) );
  AND2X1 U5942 ( .IN1(\fmul_0_0_0_0_10/sub_1_root_add_321/A[0] ), .IN2(
        \fmul_0_0_0_0_10/sub_1_root_add_321/A[1] ), .Q(n14120) );
  AND2X1 U5943 ( .IN1(n14120), .IN2(\fmul_0_0_0_0_10/sub_1_root_add_321/A[2] ), 
        .Q(n14121) );
  AND2X1 U5944 ( .IN1(n14121), .IN2(\fmul_0_0_0_0_10/sub_1_root_add_321/A[3] ), 
        .Q(n14122) );
  INVX0 U5945 ( .INP(n8803), .ZN(n14992) );
  NOR2X0 U5946 ( .IN1(n13706), .IN2(n8803), .QN(n8817) );
  INVX0 U5947 ( .INP(\fmul_0_0_0_0_10/sub_1_root_add_321/A[4] ), .ZN(n14175)
         );
  NAND2X1 U5948 ( .IN1(n13498), .IN2(n13617), .QN(n10554) );
  NAND2X1 U5949 ( .IN1(n10551), .IN2(n13618), .QN(n10549) );
  INVX0 U5950 ( .INP(n10409), .ZN(n14974) );
  INVX0 U5951 ( .INP(n11437), .ZN(n14660) );
  INVX0 U5952 ( .INP(n11218), .ZN(n14702) );
  INVX0 U5953 ( .INP(n11056), .ZN(n14755) );
  INVX0 U5954 ( .INP(n10975), .ZN(n14787) );
  INVX0 U5955 ( .INP(n11354), .ZN(n14681) );
  INVX0 U5956 ( .INP(n10732), .ZN(n14850) );
  INVX0 U5957 ( .INP(n10894), .ZN(n14808) );
  INVX0 U5958 ( .INP(n10649), .ZN(n14882) );
  INVX0 U5959 ( .INP(n10813), .ZN(n14829) );
  INVX0 U5960 ( .INP(n11137), .ZN(n14734) );
  NAND2X1 U5961 ( .IN1(n10409), .IN2(n14979), .QN(n12794) );
  INVX0 U5962 ( .INP(
        \add_0_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .ZN(n14522) );
  INVX0 U5963 ( .INP(
        \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ), .ZN(
        n14523) );
  NOR2X0 U5964 ( .IN1(\fadd_0_0_0_0_8/fracresultfar0 [6]), .IN2(
        \fadd_0_0_0_0_8/fracresultfar0 [7]), .QN(\fadd_0_0_0_0_8/add_859/B[1] ) );
  INVX0 U5965 ( .INP(n8240), .ZN(n14860) );
  NOR2X0 U5966 ( .IN1(\fadd_0_0_0_0_4/fracresultfar0 [6]), .IN2(
        \fadd_0_0_0_0_4/fracresultfar0 [7]), .QN(\fadd_0_0_0_0_4/add_859/B[1] ) );
  INVX0 U5967 ( .INP(n8407), .ZN(n14765) );
  NOR2X0 U5968 ( .IN1(\fadd_0_0_0_0_2/fracresultfar0 [6]), .IN2(
        \fadd_0_0_0_0_2/fracresultfar0 [7]), .QN(\fadd_0_0_0_0_2/add_859/B[1] ) );
  XNOR2X1 U5969 ( .IN1(
        \add_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [9]), .IN2(\fadd_0_0_0_0_8/resultbeforeround [9]), .Q(n14123) );
  INVX0 U5970 ( .INP(n8245), .ZN(n14858) );
  XNOR2X1 U5971 ( .IN1(
        \add_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [9]), .IN2(\fadd_0_0_0_0_4/resultbeforeround [9]), .Q(n14124) );
  INVX0 U5972 ( .INP(n10719), .ZN(n14849) );
  INVX0 U5973 ( .INP(n11424), .ZN(n14659) );
  INVX0 U5974 ( .INP(n10881), .ZN(n14807) );
  INVX0 U5975 ( .INP(n11205), .ZN(n14701) );
  INVX0 U5976 ( .INP(n10636), .ZN(n14881) );
  INVX0 U5977 ( .INP(n11043), .ZN(n14754) );
  INVX0 U5978 ( .INP(n10800), .ZN(n14828) );
  INVX0 U5979 ( .INP(n10962), .ZN(n14786) );
  INVX0 U5980 ( .INP(n11124), .ZN(n14733) );
  INVX0 U5981 ( .INP(n11341), .ZN(n14680) );
  XNOR2X1 U5982 ( .IN1(
        \add_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [9]), .IN2(\fadd_0_0_0_0_2/resultbeforeround [9]), .Q(n14125) );
  INVX0 U5983 ( .INP(n8996), .ZN(n14763) );
  INVX0 U5984 ( .INP(n8998), .ZN(n14710) );
  INVX0 U5985 ( .INP(\fmul_0_0_0_0_10/add_2_root_add_321/carry[5] ), .ZN(
        n14173) );
  NAND2X1 U5986 ( .IN1(n10719), .IN2(n14853), .QN(
        \fadd_0_0_0_0_8/fracyclose1 [4]) );
  NAND2X1 U5987 ( .IN1(n10636), .IN2(n14885), .QN(
        \fadd_0_0_0_0_9/fracyclose1 [4]) );
  NAND2X1 U5988 ( .IN1(n11424), .IN2(n14663), .QN(
        \fadd_0_0_0_0_0/fracyclose1 [4]) );
  NAND2X1 U5989 ( .IN1(n11043), .IN2(n14758), .QN(
        \fadd_0_0_0_0_4/fracyclose1 [4]) );
  NAND2X1 U5990 ( .IN1(n10881), .IN2(n14811), .QN(
        \fadd_0_0_0_0_6/fracyclose1 [4]) );
  NAND2X1 U5991 ( .IN1(n10800), .IN2(n14832), .QN(
        \fadd_0_0_0_0_7/fracyclose1 [4]) );
  NAND2X1 U5992 ( .IN1(n10962), .IN2(n14790), .QN(
        \fadd_0_0_0_0_5/fracyclose1 [4]) );
  NAND2X1 U5993 ( .IN1(n11124), .IN2(n14737), .QN(
        \fadd_0_0_0_0_3/fracyclose1 [4]) );
  NAND2X1 U5994 ( .IN1(n11205), .IN2(n14705), .QN(
        \fadd_0_0_0_0_2/fracyclose1 [4]) );
  NAND2X1 U5995 ( .IN1(n11341), .IN2(n14684), .QN(
        \fadd_0_0_0_0_1/fracyclose1 [4]) );
  NAND2X1 U5996 ( .IN1(n13468), .IN2(n13499), .QN(n10539) );
  INVX0 U5997 ( .INP(
        \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/n297_o[3] ), .ZN(
        n14524) );
  INVX0 U5998 ( .INP(n8219), .ZN(n14861) );
  INVX0 U5999 ( .INP(n8557), .ZN(n14713) );
  NAND2X1 U6000 ( .IN1(n13499), .IN2(n13619), .QN(n10534) );
  NOR2X0 U6001 ( .IN1(\fadd_0_0_0_0_0/fracresultfar0 [6]), .IN2(
        \fadd_0_0_0_0_0/fracresultfar0 [7]), .QN(\fadd_0_0_0_0_0/add_859/B[1] ) );
  NOR2X0 U6002 ( .IN1(\fadd_0_0_0_0_6/fracresultfar0 [6]), .IN2(
        \fadd_0_0_0_0_6/fracresultfar0 [7]), .QN(\fadd_0_0_0_0_6/add_859/B[1] ) );
  NOR2X0 U6003 ( .IN1(\fadd_0_0_0_0_7/fracresultfar0 [6]), .IN2(
        \fadd_0_0_0_0_7/fracresultfar0 [7]), .QN(\fadd_0_0_0_0_7/add_859/B[1] ) );
  NOR2X0 U6004 ( .IN1(\fadd_0_0_0_0_5/fracresultfar0 [6]), .IN2(
        \fadd_0_0_0_0_5/fracresultfar0 [7]), .QN(\fadd_0_0_0_0_5/add_859/B[1] ) );
  NOR2X0 U6005 ( .IN1(\fadd_0_0_0_0_9/fracresultfar0 [6]), .IN2(
        \fadd_0_0_0_0_9/fracresultfar0 [7]), .QN(\fadd_0_0_0_0_9/add_859/B[1] ) );
  NOR2X0 U6006 ( .IN1(\fadd_0_0_0_0_3/fracresultfar0 [6]), .IN2(
        \fadd_0_0_0_0_3/fracresultfar0 [7]), .QN(\fadd_0_0_0_0_3/add_859/B[1] ) );
  NOR2X0 U6007 ( .IN1(\fadd_0_0_0_0_1/fracresultfar0 [6]), .IN2(
        \fadd_0_0_0_0_1/fracresultfar0 [7]), .QN(\fadd_0_0_0_0_1/add_859/B[1] ) );
  INVX0 U6008 ( .INP(n8222), .ZN(n14862) );
  INVX0 U6009 ( .INP(n8527), .ZN(n14714) );
  INVX0 U6010 ( .INP(n8225), .ZN(n14863) );
  INVX0 U6011 ( .INP(n8530), .ZN(n14715) );
  INVX0 U6012 ( .INP(\fmul_0_0_0_0_10/roundingadder/add_1_root_add_57/SUM[10] ), .ZN(n14961) );
  NAND2X1 U6013 ( .IN1(n10540), .IN2(n13620), .QN(n10521) );
  INVX0 U6014 ( .INP(n10509), .ZN(n14921) );
  INVX0 U6015 ( .INP(n8228), .ZN(n14864) );
  INVX0 U6016 ( .INP(n8533), .ZN(n14716) );
  INVX0 U6017 ( .INP(
        \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ), .ZN(
        n14525) );
  INVX0 U6018 ( .INP(n8231), .ZN(n14865) );
  INVX0 U6019 ( .INP(n8536), .ZN(n14717) );
  NAND2X1 U6020 ( .IN1(\fadd_0_0_0_0_8/fracresultfar0 [6]), .IN2(n14871), .QN(
        \fadd_0_0_0_0_8/expoperationsel[0] ) );
  INVX0 U6021 ( .INP(\fadd_0_0_0_0_8/fracresultfar0 [7]), .ZN(n14871) );
  NAND2X1 U6022 ( .IN1(\fadd_0_0_0_0_4/fracresultfar0 [6]), .IN2(n14776), .QN(
        \fadd_0_0_0_0_4/expoperationsel[0] ) );
  INVX0 U6023 ( .INP(\fadd_0_0_0_0_4/fracresultfar0 [7]), .ZN(n14776) );
  NAND2X1 U6024 ( .IN1(\fadd_0_0_0_0_2/fracresultfar0 [6]), .IN2(n14723), .QN(
        \fadd_0_0_0_0_2/expoperationsel[0] ) );
  INVX0 U6025 ( .INP(\fadd_0_0_0_0_2/fracresultfar0 [7]), .ZN(n14723) );
  INVX0 U6026 ( .INP(n10692), .ZN(n14848) );
  INVX0 U6027 ( .INP(n10856), .ZN(n14806) );
  INVX0 U6028 ( .INP(n10611), .ZN(n14880) );
  INVX0 U6029 ( .INP(n10775), .ZN(n14827) );
  INVX0 U6030 ( .INP(n11099), .ZN(n14732) );
  INVX0 U6031 ( .INP(n8234), .ZN(n14866) );
  INVX0 U6032 ( .INP(n11397), .ZN(n14658) );
  INVX0 U6033 ( .INP(n11180), .ZN(n14700) );
  INVX0 U6034 ( .INP(n11018), .ZN(n14753) );
  INVX0 U6035 ( .INP(n10937), .ZN(n14785) );
  INVX0 U6036 ( .INP(n11316), .ZN(n14679) );
  INVX0 U6037 ( .INP(n8539), .ZN(n14718) );
  INVX0 U6038 ( .INP(n8237), .ZN(n14867) );
  INVX0 U6039 ( .INP(n8542), .ZN(n14719) );
  NOR2X0 U6040 ( .IN1(n10719), .IN2(n10715), .QN(n10717) );
  NOR2X0 U6041 ( .IN1(n10636), .IN2(n10632), .QN(n10634) );
  NOR2X0 U6042 ( .IN1(n10800), .IN2(n10796), .QN(n10798) );
  NOR2X0 U6043 ( .IN1(n11424), .IN2(n11420), .QN(n11422) );
  NOR2X0 U6044 ( .IN1(n11043), .IN2(n11039), .QN(n11041) );
  NOR2X0 U6045 ( .IN1(n10881), .IN2(n10877), .QN(n10879) );
  NOR2X0 U6046 ( .IN1(n10962), .IN2(n10958), .QN(n10960) );
  NOR2X0 U6047 ( .IN1(n11124), .IN2(n11120), .QN(n11122) );
  NOR2X0 U6048 ( .IN1(n11205), .IN2(n11201), .QN(n11203) );
  NOR2X0 U6049 ( .IN1(n11341), .IN2(n11337), .QN(n11339) );
  INVX0 U6050 ( .INP(n10404), .ZN(n14905) );
  INVX0 U6051 ( .INP(n8216), .ZN(n14868) );
  INVX0 U6052 ( .INP(n8545), .ZN(n14720) );
  NOR2X0 U6053 ( .IN1(n14842), .IN2(n14852), .QN(n10733) );
  NOR2X0 U6054 ( .IN1(n14652), .IN2(n14662), .QN(n11438) );
  NOR2X0 U6055 ( .IN1(n14800), .IN2(n14810), .QN(n10895) );
  NOR2X0 U6056 ( .IN1(n14694), .IN2(n14704), .QN(n11219) );
  NOR2X0 U6057 ( .IN1(n14874), .IN2(n14884), .QN(n10650) );
  NOR2X0 U6058 ( .IN1(n14821), .IN2(n14831), .QN(n10814) );
  NOR2X0 U6059 ( .IN1(n14747), .IN2(n14757), .QN(n11057) );
  NOR2X0 U6060 ( .IN1(n14779), .IN2(n14789), .QN(n10976) );
  NOR2X0 U6061 ( .IN1(n14726), .IN2(n14736), .QN(n11138) );
  NOR2X0 U6062 ( .IN1(n14673), .IN2(n14683), .QN(n11355) );
  INVX0 U6063 ( .INP(n8208), .ZN(n14869) );
  INVX0 U6064 ( .INP(n8548), .ZN(n14721) );
  NAND2X1 U6065 ( .IN1(\fadd_0_0_0_0_0/fracresultfar0 [6]), .IN2(n14670), .QN(
        \fadd_0_0_0_0_0/expoperationsel[0] ) );
  INVX0 U6066 ( .INP(\fadd_0_0_0_0_0/fracresultfar0 [7]), .ZN(n14670) );
  NAND2X1 U6067 ( .IN1(\fadd_0_0_0_0_6/fracresultfar0 [6]), .IN2(n14818), .QN(
        \fadd_0_0_0_0_6/expoperationsel[0] ) );
  INVX0 U6068 ( .INP(\fadd_0_0_0_0_6/fracresultfar0 [7]), .ZN(n14818) );
  NAND2X1 U6069 ( .IN1(\fadd_0_0_0_0_7/fracresultfar0 [6]), .IN2(n14839), .QN(
        \fadd_0_0_0_0_7/expoperationsel[0] ) );
  INVX0 U6070 ( .INP(\fadd_0_0_0_0_7/fracresultfar0 [7]), .ZN(n14839) );
  NAND2X1 U6071 ( .IN1(\fadd_0_0_0_0_5/fracresultfar0 [6]), .IN2(n14797), .QN(
        \fadd_0_0_0_0_5/expoperationsel[0] ) );
  INVX0 U6072 ( .INP(\fadd_0_0_0_0_5/fracresultfar0 [7]), .ZN(n14797) );
  NAND2X1 U6073 ( .IN1(\fadd_0_0_0_0_9/fracresultfar0 [6]), .IN2(n14892), .QN(
        \fadd_0_0_0_0_9/expoperationsel[0] ) );
  INVX0 U6074 ( .INP(\fadd_0_0_0_0_9/fracresultfar0 [7]), .ZN(n14892) );
  NAND2X1 U6075 ( .IN1(\fadd_0_0_0_0_3/fracresultfar0 [6]), .IN2(n14744), .QN(
        \fadd_0_0_0_0_3/expoperationsel[0] ) );
  INVX0 U6076 ( .INP(\fadd_0_0_0_0_3/fracresultfar0 [7]), .ZN(n14744) );
  NAND2X1 U6077 ( .IN1(\fadd_0_0_0_0_1/fracresultfar0 [6]), .IN2(n14691), .QN(
        \fadd_0_0_0_0_1/expoperationsel[0] ) );
  INVX0 U6078 ( .INP(\fadd_0_0_0_0_1/fracresultfar0 [7]), .ZN(n14691) );
  NOR2X0 U6079 ( .IN1(n10732), .IN2(n10723), .QN(n12771) );
  NOR2X0 U6080 ( .IN1(n11437), .IN2(n11428), .QN(n12693) );
  NOR2X0 U6081 ( .IN1(n10894), .IN2(n10885), .QN(n12753) );
  NOR2X0 U6082 ( .IN1(n11218), .IN2(n11209), .QN(n12713) );
  NOR2X0 U6083 ( .IN1(n10649), .IN2(n10640), .QN(n12781) );
  NOR2X0 U6084 ( .IN1(n11056), .IN2(n11047), .QN(n12733) );
  NOR2X0 U6085 ( .IN1(n10813), .IN2(n10804), .QN(n12761) );
  NOR2X0 U6086 ( .IN1(n10975), .IN2(n10966), .QN(n12741) );
  NOR2X0 U6087 ( .IN1(n11137), .IN2(n11128), .QN(n12721) );
  NOR2X0 U6088 ( .IN1(n11354), .IN2(n11345), .QN(n12701) );
  NOR2X0 U6089 ( .IN1(n10719), .IN2(n10723), .QN(
        \fadd_0_0_0_0_8/rightshiftercomponent/level2[1] ) );
  NOR2X0 U6090 ( .IN1(n11424), .IN2(n11428), .QN(
        \fadd_0_0_0_0_0/rightshiftercomponent/level2[1] ) );
  NOR2X0 U6091 ( .IN1(n10881), .IN2(n10885), .QN(
        \fadd_0_0_0_0_6/rightshiftercomponent/level2[1] ) );
  NOR2X0 U6092 ( .IN1(n11205), .IN2(n11209), .QN(
        \fadd_0_0_0_0_2/rightshiftercomponent/level2[1] ) );
  NOR2X0 U6093 ( .IN1(n10636), .IN2(n10640), .QN(
        \fadd_0_0_0_0_9/rightshiftercomponent/level2[1] ) );
  NOR2X0 U6094 ( .IN1(n11043), .IN2(n11047), .QN(
        \fadd_0_0_0_0_4/rightshiftercomponent/level2[1] ) );
  NOR2X0 U6095 ( .IN1(n10800), .IN2(n10804), .QN(
        \fadd_0_0_0_0_7/rightshiftercomponent/level2[1] ) );
  NOR2X0 U6096 ( .IN1(n10962), .IN2(n10966), .QN(
        \fadd_0_0_0_0_5/rightshiftercomponent/level2[1] ) );
  NOR2X0 U6097 ( .IN1(n11124), .IN2(n11128), .QN(
        \fadd_0_0_0_0_3/rightshiftercomponent/level2[1] ) );
  NOR2X0 U6098 ( .IN1(n11341), .IN2(n11345), .QN(
        \fadd_0_0_0_0_1/rightshiftercomponent/level2[1] ) );
  OR4X1 U6099 ( .IN1(n14188), .IN2(n11272), .IN3(\fadd_0_0_0_0_10/U5/DATA2_1 ), 
        .IN4(\fadd_0_0_0_0_10/U5/DATA2_2 ), .Q(n11283) );
  NAND2X1 U6100 ( .IN1(n9055), .IN2(n14263), .QN(n9009) );
  AO221X1 U6101 ( .IN1(\fadd_0_0_0_0_10/U5/DATA2_2 ), .IN2(n11271), .IN3(
        \fadd_0_0_0_0_10/U5/DATA1_2 ), .IN4(n14188), .IN5(n11263), .Q(
        \fadd_0_0_0_0_10/U27/Z_2 ) );
  AO22X1 U6102 ( .IN1(n11271), .IN2(n11272), .IN3(n11273), .IN4(n14304), .Q(
        n11263) );
  NOR2X0 U6103 ( .IN1(n10409), .IN2(n14977), .QN(n11246) );
  AO221X1 U6104 ( .IN1(\fadd_0_0_0_0_10/U5/DATA2_1 ), .IN2(n11271), .IN3(
        \fadd_0_0_0_0_10/U5/DATA1_1 ), .IN4(n14188), .IN5(n11263), .Q(
        \fadd_0_0_0_0_10/U27/Z_1 ) );
  AND2X1 U6105 ( .IN1(n9055), .IN2(n8764), .Q(n8989) );
  NOR2X0 U6106 ( .IN1(n11263), .IN2(\fadd_0_0_0_0_10/U27/DATA1_0 ), .QN(n11242) );
  NBUFFX2 U6107 ( .INP(n9441), .Z(n14396) );
  NBUFFX2 U6108 ( .INP(n9441), .Z(n14395) );
  NOR2X0 U6109 ( .IN1(n14976), .IN2(n11251), .QN(
        \fadd_0_0_0_0_10/rightshiftercomponent/U6/Z_0 ) );
  NAND2X1 U6110 ( .IN1(n14976), .IN2(n11262), .QN(n11260) );
  INVX0 U6111 ( .INP(n8997), .ZN(n14910) );
  INVX0 U6112 ( .INP(\fmul_0_0_0_0_10/sub_1_root_add_321/A[0] ), .ZN(n14919)
         );
  INVX0 U6113 ( .INP(n11280), .ZN(n14940) );
  NOR2X0 U6114 ( .IN1(\fadd_0_0_0_0_8/exponentdifferencexy [3]), .IN2(
        \fadd_0_0_0_0_8/exponentdifferencexy [4]), .QN(n10697) );
  NOR2X0 U6115 ( .IN1(\fadd_0_0_0_0_9/exponentdifferencexy [3]), .IN2(
        \fadd_0_0_0_0_9/exponentdifferencexy [4]), .QN(n10616) );
  NOR2X0 U6116 ( .IN1(\fadd_0_0_0_0_7/exponentdifferencexy [3]), .IN2(
        \fadd_0_0_0_0_7/exponentdifferencexy [4]), .QN(n10780) );
  NOR2X0 U6117 ( .IN1(\fadd_0_0_0_0_0/exponentdifferencexy [3]), .IN2(
        \fadd_0_0_0_0_0/exponentdifferencexy [4]), .QN(n11402) );
  NOR2X0 U6118 ( .IN1(\fadd_0_0_0_0_4/exponentdifferencexy [3]), .IN2(
        \fadd_0_0_0_0_4/exponentdifferencexy [4]), .QN(n11023) );
  NOR2X0 U6119 ( .IN1(\fadd_0_0_0_0_6/exponentdifferencexy [3]), .IN2(
        \fadd_0_0_0_0_6/exponentdifferencexy [4]), .QN(n10861) );
  NOR2X0 U6120 ( .IN1(\fadd_0_0_0_0_5/exponentdifferencexy [3]), .IN2(
        \fadd_0_0_0_0_5/exponentdifferencexy [4]), .QN(n10942) );
  NOR2X0 U6121 ( .IN1(\fadd_0_0_0_0_3/exponentdifferencexy [3]), .IN2(
        \fadd_0_0_0_0_3/exponentdifferencexy [4]), .QN(n11104) );
  NOR2X0 U6122 ( .IN1(\fadd_0_0_0_0_2/exponentdifferencexy [3]), .IN2(
        \fadd_0_0_0_0_2/exponentdifferencexy [4]), .QN(n11185) );
  NOR2X0 U6123 ( .IN1(\fadd_0_0_0_0_1/exponentdifferencexy [3]), .IN2(
        \fadd_0_0_0_0_1/exponentdifferencexy [4]), .QN(n11321) );
  AND2X1 U6124 ( .IN1(n9129), .IN2(n14436), .Q(n9062) );
  AND2X1 U6125 ( .IN1(n9129), .IN2(n8764), .Q(n9096) );
  NBUFFX2 U6126 ( .INP(n9450), .Z(n14363) );
  NBUFFX2 U6127 ( .INP(n9450), .Z(n14362) );
  NBUFFX2 U6128 ( .INP(n9450), .Z(n14361) );
  NBUFFX2 U6129 ( .INP(n9446), .Z(n14375) );
  NBUFFX2 U6130 ( .INP(n9447), .Z(n14374) );
  NAND2X1 U6131 ( .IN1(n14177), .IN2(n13749), .QN(
        \fadd_0_0_0_0_10/sub_784/carry[4] ) );
  INVX0 U6132 ( .INP(\fadd_0_0_0_0_10/sub_784/carry[3] ), .ZN(n14177) );
  AND2X1 U6133 ( .IN1(n14176), .IN2(n13884), .Q(n14126) );
  INVX0 U6134 ( .INP(\fadd_0_0_0_0_8/sub_784/B[0] ), .ZN(n14629) );
  INVX0 U6135 ( .INP(\fadd_0_0_0_0_9/sub_784/B[0] ), .ZN(n14640) );
  INVX0 U6136 ( .INP(\fadd_0_0_0_0_0/sub_784/B[0] ), .ZN(n14541) );
  INVX0 U6137 ( .INP(\fadd_0_0_0_0_4/sub_784/B[0] ), .ZN(n14585) );
  INVX0 U6138 ( .INP(\fadd_0_0_0_0_6/sub_784/B[0] ), .ZN(n14607) );
  INVX0 U6139 ( .INP(\fadd_0_0_0_0_7/sub_784/B[0] ), .ZN(n14618) );
  INVX0 U6140 ( .INP(\fadd_0_0_0_0_5/sub_784/B[0] ), .ZN(n14596) );
  INVX0 U6141 ( .INP(\fadd_0_0_0_0_2/sub_784/B[0] ), .ZN(n14563) );
  INVX0 U6142 ( .INP(\fadd_0_0_0_0_3/sub_784/B[0] ), .ZN(n14574) );
  INVX0 U6143 ( .INP(\fadd_0_0_0_0_1/sub_784/B[0] ), .ZN(n14552) );
  NOR2X0 U6144 ( .IN1(n10503), .IN2(n14921), .QN(n10500) );
  INVX0 U6145 ( .INP(n10502), .ZN(n14922) );
  NAND2X1 U6146 ( .IN1(n10509), .IN2(n10510), .QN(n10506) );
  NOR2X0 U6147 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/carry [5]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/A[5] ), .QN(n14127)
         );
  INVX0 U6148 ( .INP(n10393), .ZN(n14915) );
  NOR2X0 U6149 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/carry [5]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/A[5] ), .QN(n14128)
         );
  NOR2X0 U6150 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/carry [5]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/A[5] ), .QN(n14129)
         );
  NOR2X0 U6151 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/carry [5]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/A[5] ), .QN(n14130)
         );
  NOR2X0 U6152 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/carry [5]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/A[5] ), .QN(n14131)
         );
  NOR2X0 U6153 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/carry [5]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/A[5] ), .QN(n14132)
         );
  NOR2X0 U6154 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/carry [5]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/A[5] ), .QN(n14133)
         );
  NOR2X0 U6155 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/carry [5]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/A[5] ), .QN(n14134)
         );
  NOR2X0 U6156 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/carry [5]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/A[5] ), .QN(n14135)
         );
  NOR2X0 U6157 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/carry [5]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/A[5] ), .QN(n14136)
         );
  INVX0 U6158 ( .INP(n14282), .ZN(n14281) );
  INVX0 U6159 ( .INP(n14301), .ZN(n14300) );
  NBUFFX2 U6160 ( .INP(n9454), .Z(n14324) );
  INVX0 U6161 ( .INP(\fadd_0_0_0_0_8/exponentdifferencexy [2]), .ZN(n14854) );
  INVX0 U6162 ( .INP(\fadd_0_0_0_0_9/exponentdifferencexy [2]), .ZN(n14886) );
  INVX0 U6163 ( .INP(\fadd_0_0_0_0_7/exponentdifferencexy [2]), .ZN(n14833) );
  INVX0 U6164 ( .INP(\fadd_0_0_0_0_0/exponentdifferencexy [2]), .ZN(n14664) );
  INVX0 U6165 ( .INP(\fadd_0_0_0_0_4/exponentdifferencexy [2]), .ZN(n14759) );
  INVX0 U6166 ( .INP(\fadd_0_0_0_0_6/exponentdifferencexy [2]), .ZN(n14812) );
  INVX0 U6167 ( .INP(\fadd_0_0_0_0_5/exponentdifferencexy [2]), .ZN(n14791) );
  INVX0 U6168 ( .INP(\fadd_0_0_0_0_3/exponentdifferencexy [2]), .ZN(n14738) );
  INVX0 U6169 ( .INP(\fadd_0_0_0_0_2/exponentdifferencexy [2]), .ZN(n14706) );
  INVX0 U6170 ( .INP(\fadd_0_0_0_0_1/exponentdifferencexy [2]), .ZN(n14685) );
  INVX0 U6171 ( .INP(\fadd_0_0_0_0_8/exponentdifferenceyx [2]), .ZN(n14856) );
  INVX0 U6172 ( .INP(\fadd_0_0_0_0_9/exponentdifferenceyx [2]), .ZN(n14888) );
  INVX0 U6173 ( .INP(\fadd_0_0_0_0_7/exponentdifferenceyx [2]), .ZN(n14835) );
  INVX0 U6174 ( .INP(\fadd_0_0_0_0_0/exponentdifferenceyx [2]), .ZN(n14666) );
  INVX0 U6175 ( .INP(\fadd_0_0_0_0_4/exponentdifferenceyx [2]), .ZN(n14761) );
  INVX0 U6176 ( .INP(\fadd_0_0_0_0_6/exponentdifferenceyx [2]), .ZN(n14814) );
  INVX0 U6177 ( .INP(\fadd_0_0_0_0_5/exponentdifferenceyx [2]), .ZN(n14793) );
  INVX0 U6178 ( .INP(\fadd_0_0_0_0_3/exponentdifferenceyx [2]), .ZN(n14740) );
  INVX0 U6179 ( .INP(\fadd_0_0_0_0_2/exponentdifferenceyx [2]), .ZN(n14708) );
  INVX0 U6180 ( .INP(\fadd_0_0_0_0_1/exponentdifferenceyx [2]), .ZN(n14687) );
  NBUFFX2 U6181 ( .INP(n9455), .Z(n14323) );
  INVX0 U6182 ( .INP(n8732), .ZN(n14918) );
  INVX0 U6183 ( .INP(\fadd_0_0_0_0_8/exponentdifferencexy [1]), .ZN(n14855) );
  INVX0 U6184 ( .INP(\fadd_0_0_0_0_9/exponentdifferencexy [1]), .ZN(n14887) );
  INVX0 U6185 ( .INP(\fadd_0_0_0_0_7/exponentdifferencexy [1]), .ZN(n14834) );
  INVX0 U6186 ( .INP(\fadd_0_0_0_0_0/exponentdifferencexy [1]), .ZN(n14665) );
  INVX0 U6187 ( .INP(\fadd_0_0_0_0_4/exponentdifferencexy [1]), .ZN(n14760) );
  INVX0 U6188 ( .INP(\fadd_0_0_0_0_6/exponentdifferencexy [1]), .ZN(n14813) );
  INVX0 U6189 ( .INP(\fadd_0_0_0_0_5/exponentdifferencexy [1]), .ZN(n14792) );
  INVX0 U6190 ( .INP(\fadd_0_0_0_0_3/exponentdifferencexy [1]), .ZN(n14739) );
  INVX0 U6191 ( .INP(\fadd_0_0_0_0_2/exponentdifferencexy [1]), .ZN(n14707) );
  INVX0 U6192 ( .INP(\fadd_0_0_0_0_1/exponentdifferencexy [1]), .ZN(n14686) );
  INVX0 U6193 ( .INP(\fadd_0_0_0_0_8/exponentdifferenceyx [1]), .ZN(n14857) );
  INVX0 U6194 ( .INP(\fadd_0_0_0_0_9/exponentdifferenceyx [1]), .ZN(n14889) );
  INVX0 U6195 ( .INP(\fadd_0_0_0_0_7/exponentdifferenceyx [1]), .ZN(n14836) );
  INVX0 U6196 ( .INP(\fadd_0_0_0_0_0/exponentdifferenceyx [1]), .ZN(n14667) );
  INVX0 U6197 ( .INP(\fadd_0_0_0_0_4/exponentdifferenceyx [1]), .ZN(n14762) );
  INVX0 U6198 ( .INP(\fadd_0_0_0_0_6/exponentdifferenceyx [1]), .ZN(n14815) );
  INVX0 U6199 ( .INP(\fadd_0_0_0_0_5/exponentdifferenceyx [1]), .ZN(n14794) );
  INVX0 U6200 ( .INP(\fadd_0_0_0_0_3/exponentdifferenceyx [1]), .ZN(n14741) );
  INVX0 U6201 ( .INP(\fadd_0_0_0_0_2/exponentdifferenceyx [1]), .ZN(n14709) );
  INVX0 U6202 ( .INP(\fadd_0_0_0_0_1/exponentdifferenceyx [1]), .ZN(n14688) );
  INVX0 U6203 ( .INP(\fmul_0_0_0_0_4/expsigpostround [10]), .ZN(n14898) );
  NOR2X0 U6204 ( .IN1(n10576), .IN2(n10577), .QN(\fmul_0_0_0_0_0/round ) );
  NOR4X0 U6205 ( .IN1(n10578), .IN2(\fmul_0_0_0_0_0/sigprod [0]), .IN3(
        \fmul_0_0_0_0_0/sigprod [2]), .IN4(\fmul_0_0_0_0_0/sigprod [1]), .QN(
        n10576) );
  INVX0 U6206 ( .INP(\fmul_0_0_0_0_3/expsigpostround [10]), .ZN(n14897) );
  INVX0 U6207 ( .INP(\fmul_0_0_0_0_1/expsigpostround [10]), .ZN(n14895) );
  INVX0 U6208 ( .INP(\fmul_0_0_0_0_5/expsigpostround [10]), .ZN(n14899) );
  INVX0 U6209 ( .INP(\fmul_0_0_0_0_7/expsigpostround [10]), .ZN(n14901) );
  INVX0 U6210 ( .INP(\fmul_0_0_0_0_2/expsigpostround [10]), .ZN(n14896) );
  INVX0 U6211 ( .INP(\fmul_0_0_0_0_9/expsigpostround [10]), .ZN(n14903) );
  INVX0 U6212 ( .INP(\fmul_0_0_0_0_6/expsigpostround [10]), .ZN(n14900) );
  NBUFFX2 U6213 ( .INP(n14200), .Z(n14258) );
  NAND2X1 U6214 ( .IN1(n10419), .IN2(n14937), .QN(n10626) );
  NAND2X1 U6215 ( .IN1(n10418), .IN2(n14936), .QN(n10707) );
  NAND2X1 U6216 ( .IN1(n10417), .IN2(n14935), .QN(n10790) );
  NAND2X1 U6217 ( .IN1(n10416), .IN2(n14934), .QN(n10871) );
  NAND2X1 U6218 ( .IN1(n10415), .IN2(n14933), .QN(n10952) );
  NAND2X1 U6219 ( .IN1(n10414), .IN2(n14932), .QN(n11033) );
  NAND2X1 U6220 ( .IN1(n10413), .IN2(n14931), .QN(n11114) );
  NAND2X1 U6221 ( .IN1(n10412), .IN2(n14930), .QN(n11195) );
  NAND2X1 U6222 ( .IN1(n10411), .IN2(n14929), .QN(n11331) );
  NAND2X1 U6223 ( .IN1(n10410), .IN2(n14928), .QN(n11412) );
  INVX0 U6224 ( .INP(n8683), .ZN(n15001) );
  INVX0 U6225 ( .INP(n9068), .ZN(n14955) );
  INVX0 U6226 ( .INP(n9288), .ZN(n14945) );
  INVX0 U6227 ( .INP(n8774), .ZN(n14986) );
  INVX0 U6228 ( .INP(n9010), .ZN(n14954) );
  NAND2X1 U6229 ( .IN1(n12870), .IN2(n12871), .QN(n11238) );
  INVX0 U6230 ( .INP(n8523), .ZN(n14944) );
  INVX0 U6231 ( .INP(n9139), .ZN(n14952) );
  INVX0 U6232 ( .INP(n8910), .ZN(n14959) );
  INVX0 U6233 ( .INP(n9350), .ZN(n14943) );
  INVX0 U6234 ( .INP(n9392), .ZN(n14941) );
  INVX0 U6235 ( .INP(n8958), .ZN(n14957) );
  INVX0 U6236 ( .INP(n9202), .ZN(n14950) );
  INVX0 U6237 ( .INP(n9244), .ZN(n14948) );
  NBUFFX2 U6238 ( .INP(n14916), .Z(n14260) );
  NBUFFX2 U6239 ( .INP(n14916), .Z(n14261) );
  NBUFFX2 U6240 ( .INP(n14916), .Z(n14259) );
  NBUFFX2 U6241 ( .INP(n14916), .Z(n14262) );
  NAND2X1 U6242 ( .IN1(n8766), .IN2(n12828), .QN(n9130) );
  NAND3X0 U6243 ( .IN1(n12826), .IN2(n14251), .IN3(n11959), .QN(n8680) );
  NAND2X1 U6244 ( .IN1(n8709), .IN2(n8710), .QN(n12883) );
  NAND2X1 U6245 ( .IN1(n8707), .IN2(n8708), .QN(n12882) );
  NAND2X1 U6246 ( .IN1(n8693), .IN2(n8694), .QN(n12875) );
  NAND2X1 U6247 ( .IN1(n8695), .IN2(n8696), .QN(n12876) );
  NAND2X1 U6248 ( .IN1(n8697), .IN2(n8698), .QN(n12877) );
  NAND2X1 U6249 ( .IN1(n8699), .IN2(n8700), .QN(n12878) );
  NAND2X1 U6250 ( .IN1(n8701), .IN2(n8702), .QN(n12879) );
  NAND2X1 U6251 ( .IN1(n8703), .IN2(n8704), .QN(n12880) );
  NAND2X1 U6252 ( .IN1(n8705), .IN2(n8706), .QN(n12881) );
  NAND2X1 U6253 ( .IN1(n8681), .IN2(n8682), .QN(n12873) );
  NAND2X1 U6254 ( .IN1(n8671), .IN2(n8672), .QN(n12872) );
  NAND2X1 U6255 ( .IN1(n8686), .IN2(n8687), .QN(n12874) );
  NAND2X1 U6256 ( .IN1(n8723), .IN2(n8724), .QN(n12885) );
  NAND2X1 U6257 ( .IN1(n8726), .IN2(n13753), .QN(n8725) );
  NAND2X1 U6258 ( .IN1(n8713), .IN2(n8714), .QN(n12884) );
  NOR2X0 U6259 ( .IN1(n8717), .IN2(n11961), .QN(n8715) );
  NAND2X1 U6260 ( .IN1(n8730), .IN2(n8731), .QN(n12886) );
  INVX0 U6261 ( .INP(\U120/DATA1_9 ), .ZN(n14904) );
  NAND2X1 U6262 ( .IN1(n13780), .IN2(n9171), .QN(n9167) );
  NOR2X0 U6263 ( .IN1(\fmul_0_0_0_0_6/expsigpostround [9]), .IN2(
        \fmul_0_0_0_0_6/expsigpostround [10]), .QN(n9177) );
  NOR2X0 U6264 ( .IN1(n13736), .IN2(n12830), .QN(n9440) );
  AO221X1 U6265 ( .IN1(n9441), .IN2(n10391), .IN3(\U571/DATA1_0 ), .IN4(n13736), .IN5(n10392), .Q(n9436) );
  AO21X1 U6266 ( .IN1(n5954), .IN2(n14242), .IN3(n9436), .Q(n13399) );
  AO21X1 U6267 ( .IN1(n5882), .IN2(n14245), .IN3(n9436), .Q(n13352) );
  AO21X1 U6268 ( .IN1(n5810), .IN2(n14234), .IN3(n9436), .Q(n13328) );
  AO21X1 U6269 ( .IN1(n5738), .IN2(n14246), .IN3(n9436), .Q(n13304) );
  AO21X1 U6270 ( .IN1(n5666), .IN2(n14246), .IN3(n9436), .Q(n13280) );
  AO21X1 U6271 ( .IN1(n5594), .IN2(n14242), .IN3(n9436), .Q(n13256) );
  AO21X1 U6272 ( .IN1(n5522), .IN2(n14242), .IN3(n9436), .Q(n13232) );
  AO21X1 U6273 ( .IN1(n5450), .IN2(n14243), .IN3(n9436), .Q(n13208) );
  AO21X1 U6274 ( .IN1(n5378), .IN2(n14243), .IN3(n9436), .Q(n13184) );
  AO21X1 U6275 ( .IN1(n5306), .IN2(n14244), .IN3(n9436), .Q(n13160) );
  NAND2X1 U6276 ( .IN1(n13781), .IN2(n9319), .QN(n9315) );
  NOR2X0 U6277 ( .IN1(\fmul_0_0_0_0_2/expsigpostround [9]), .IN2(
        \fmul_0_0_0_0_2/expsigpostround [10]), .QN(n9325) );
  AO221X1 U6278 ( .IN1(n14395), .IN2(n10385), .IN3(\U576/DATA1_1 ), .IN4(n9440), .IN5(n10386), .Q(n9544) );
  AO221X1 U6279 ( .IN1(n14396), .IN2(n10379), .IN3(\U576/DATA1_2 ), .IN4(n9440), .IN5(n10380), .Q(n9542) );
  AO221X1 U6280 ( .IN1(n9441), .IN2(n10373), .IN3(\U576/DATA1_3 ), .IN4(n9440), 
        .IN5(n10374), .Q(n9540) );
  AO221X1 U6281 ( .IN1(n9441), .IN2(n10367), .IN3(\U576/DATA1_4 ), .IN4(n9440), 
        .IN5(n10368), .Q(n9538) );
  AO221X1 U6282 ( .IN1(n9441), .IN2(n10361), .IN3(\U576/DATA1_5 ), .IN4(n9440), 
        .IN5(n10362), .Q(n9537) );
  AO221X1 U6283 ( .IN1(n9441), .IN2(n10355), .IN3(\U576/DATA1_6 ), .IN4(n9440), 
        .IN5(n10356), .Q(n9536) );
  AO221X1 U6284 ( .IN1(n9441), .IN2(n10349), .IN3(\U576/DATA1_7 ), .IN4(n9440), 
        .IN5(n10350), .Q(n9535) );
  AO221X1 U6285 ( .IN1(n14396), .IN2(n10343), .IN3(\U576/DATA1_8 ), .IN4(n9440), .IN5(n10344), .Q(n9534) );
  AO221X1 U6286 ( .IN1(n9441), .IN2(n10337), .IN3(\U576/DATA1_9 ), .IN4(n9440), 
        .IN5(n10338), .Q(n9533) );
  AO221X1 U6287 ( .IN1(n9441), .IN2(n10330), .IN3(\U576/DATA1_10 ), .IN4(n9440), .IN5(n10331), .Q(n9531) );
  AO221X1 U6288 ( .IN1(n9441), .IN2(n10323), .IN3(\U576/DATA1_11 ), .IN4(
        n14406), .IN5(n10324), .Q(n9529) );
  NOR2X0 U6289 ( .IN1(n14437), .IN2(n12143), .QN(\U4/Z_50 ) );
  NOR2X0 U6290 ( .IN1(n14437), .IN2(n12009), .QN(\U4/Z_49 ) );
  NOR2X0 U6291 ( .IN1(n14437), .IN2(n12826), .QN(\U4/Z_46 ) );
  NOR2X0 U6292 ( .IN1(rst), .IN2(n11468), .QN(\U4/Z_53 ) );
  NOR2X0 U6293 ( .IN1(n14437), .IN2(n11466), .QN(\U4/Z_48 ) );
  NOR2X0 U6294 ( .IN1(n14437), .IN2(n11464), .QN(\U4/Z_43 ) );
  NOR2X0 U6295 ( .IN1(n14437), .IN2(n11952), .QN(\U4/Z_47 ) );
  NOR2X0 U6296 ( .IN1(n14437), .IN2(n11959), .QN(\U4/Z_51 ) );
  NOR2X0 U6297 ( .IN1(rst), .IN2(n12007), .QN(\U4/Z_54 ) );
  NOR2X0 U6298 ( .IN1(rst), .IN2(n12836), .QN(n13436) );
  NOR2X0 U6299 ( .IN1(rst), .IN2(n12837), .QN(n13439) );
  NOR2X0 U6300 ( .IN1(rst), .IN2(n11937), .QN(n13440) );
  NOR2X0 U6301 ( .IN1(rst), .IN2(n11467), .QN(\U4/Z_52 ) );
  NOR2X0 U6302 ( .IN1(n14437), .IN2(n11465), .QN(\U4/Z_45 ) );
  NOR2X0 U6303 ( .IN1(n14437), .IN2(n11463), .QN(\U4/Z_42 ) );
  NOR2X0 U6304 ( .IN1(rst), .IN2(n11611), .QN(n13435) );
  NOR2X0 U6305 ( .IN1(rst), .IN2(n11610), .QN(n13438) );
  NOR2X0 U6306 ( .IN1(rst), .IN2(n11608), .QN(n13441) );
  NOR2X0 U6307 ( .IN1(n14437), .IN2(n12828), .QN(\U4/Z_41 ) );
  OR2X1 U6308 ( .IN1(n14187), .IN2(n12829), .Q(n14137) );
  NOR2X0 U6309 ( .IN1(n14439), .IN2(n12833), .QN(\U4/Z_16 ) );
  NOR2X0 U6310 ( .IN1(n14439), .IN2(n12832), .QN(\U4/Z_19 ) );
  NOR2X0 U6311 ( .IN1(n14438), .IN2(n12830), .QN(\U4/Z_28 ) );
  NOR2X0 U6312 ( .IN1(n14439), .IN2(n12831), .QN(\U4/Z_25 ) );
  NOR2X0 U6313 ( .IN1(n14438), .IN2(n11928), .QN(\U4/Z_31 ) );
  NOR2X0 U6314 ( .IN1(n14439), .IN2(n11930), .QN(\U4/Z_15 ) );
  NOR2X0 U6315 ( .IN1(n14439), .IN2(n11931), .QN(\U4/Z_18 ) );
  NOR2X0 U6316 ( .IN1(n14439), .IN2(n11932), .QN(\U4/Z_21 ) );
  NOR2X0 U6317 ( .IN1(n14438), .IN2(n11934), .QN(\U4/Z_27 ) );
  NOR2X0 U6318 ( .IN1(n14439), .IN2(n11933), .QN(\U4/Z_24 ) );
  NOR2X0 U6319 ( .IN1(n14438), .IN2(n11462), .QN(\U4/Z_39 ) );
  NOR2X0 U6320 ( .IN1(n14438), .IN2(n11461), .QN(\U4/Z_38 ) );
  NOR2X0 U6321 ( .IN1(n14438), .IN2(n11460), .QN(\U4/Z_35 ) );
  NOR2X0 U6322 ( .IN1(n14438), .IN2(n11459), .QN(\U4/Z_34 ) );
  NOR2X0 U6323 ( .IN1(n14438), .IN2(n11458), .QN(\U4/Z_32 ) );
  NOR2X0 U6324 ( .IN1(n14438), .IN2(n11457), .QN(\U4/Z_29 ) );
  NOR2X0 U6325 ( .IN1(n14438), .IN2(n11456), .QN(\U4/Z_26 ) );
  NOR2X0 U6326 ( .IN1(n14439), .IN2(n11455), .QN(\U4/Z_23 ) );
  NOR2X0 U6327 ( .IN1(n14439), .IN2(n11454), .QN(\U4/Z_20 ) );
  NOR2X0 U6328 ( .IN1(n14439), .IN2(n11453), .QN(\U4/Z_17 ) );
  NOR2X0 U6329 ( .IN1(n14439), .IN2(n11452), .QN(\U4/Z_14 ) );
  NOR2X0 U6330 ( .IN1(n14439), .IN2(n12835), .QN(\U4/Z_10 ) );
  NOR2X0 U6331 ( .IN1(n14438), .IN2(n12834), .QN(\U4/Z_13 ) );
  NOR2X0 U6332 ( .IN1(n14439), .IN2(n11929), .QN(\U4/Z_12 ) );
  NOR2X0 U6333 ( .IN1(n14438), .IN2(n11451), .QN(\U4/Z_11 ) );
  NAND2X1 U6334 ( .IN1(n13750), .IN2(n9102), .QN(n9100) );
  NOR2X0 U6335 ( .IN1(\fmul_0_0_0_0_4/expsigpostround [9]), .IN2(
        \fmul_0_0_0_0_4/expsigpostround [10]), .QN(n9108) );
  AND3X1 U6336 ( .IN1(n12827), .IN2(n8997), .IN3(n11952), .Q(n9055) );
  OR2X1 U6337 ( .IN1(n14162), .IN2(n14419), .Q(n8997) );
  NAND2X1 U6338 ( .IN1(n9011), .IN2(n9012), .QN(n12959) );
  INVX0 U6339 ( .INP(n8380), .ZN(n14766) );
  NAND2X1 U6340 ( .IN1(n9016), .IN2(n9017), .QN(n12960) );
  INVX0 U6341 ( .INP(n8383), .ZN(n14767) );
  NAND2X1 U6342 ( .IN1(n9021), .IN2(n9022), .QN(n12961) );
  INVX0 U6343 ( .INP(n8386), .ZN(n14768) );
  NAND2X1 U6344 ( .IN1(n9026), .IN2(n9027), .QN(n12962) );
  INVX0 U6345 ( .INP(n8389), .ZN(n14769) );
  NAND2X1 U6346 ( .IN1(n9031), .IN2(n9032), .QN(n12963) );
  INVX0 U6347 ( .INP(n8392), .ZN(n14770) );
  NAND2X1 U6348 ( .IN1(n9036), .IN2(n9037), .QN(n12964) );
  INVX0 U6349 ( .INP(n8395), .ZN(n14771) );
  NAND2X1 U6350 ( .IN1(n9041), .IN2(n9042), .QN(n12965) );
  INVX0 U6351 ( .INP(n8398), .ZN(n14772) );
  NAND2X1 U6352 ( .IN1(n9046), .IN2(n9047), .QN(n12966) );
  INVX0 U6353 ( .INP(n8401), .ZN(n14773) );
  NAND2X1 U6354 ( .IN1(n9051), .IN2(n9052), .QN(n12967) );
  INVX0 U6355 ( .INP(n8404), .ZN(n14774) );
  NAND2X1 U6356 ( .IN1(n9007), .IN2(n9008), .QN(n12958) );
  NAND2X1 U6357 ( .IN1(n9000), .IN2(n9001), .QN(n12957) );
  INVX0 U6358 ( .INP(n8551), .ZN(n14712) );
  NAND2X1 U6359 ( .IN1(n8991), .IN2(n8992), .QN(n12956) );
  NAND2X1 U6360 ( .IN1(n11953), .IN2(n8994), .QN(n8993) );
  NAND2X1 U6361 ( .IN1(n8777), .IN2(n8778), .QN(n8781) );
  NAND2X1 U6362 ( .IN1(n13632), .IN2(n14171), .QN(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/carry[7] ) );
  NOR4X0 U6363 ( .IN1(n12070), .IN2(n12071), .IN3(n12072), .IN4(n12073), .QN(
        n8776) );
  INVX0 U6364 ( .INP(n8770), .ZN(n14984) );
  AND2X1 U6365 ( .IN1(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/B[1] ), .IN2(n14139), .Q(n14138) );
  NOR2X0 U6366 ( .IN1(n12062), .IN2(n12063), .QN(n8879) );
  AND2X1 U6367 ( .IN1(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/B[0] ), .IN2(\fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/CI ), 
        .Q(n14139) );
  NAND2X1 U6368 ( .IN1(n8869), .IN2(n12068), .QN(n8838) );
  NAND2X1 U6369 ( .IN1(n12068), .IN2(n13412), .QN(n8805) );
  NAND2X1 U6370 ( .IN1(n8791), .IN2(n8790), .QN(n8799) );
  NAND2X1 U6371 ( .IN1(n13885), .IN2(n14180), .QN(
        \fadd_0_0_0_0_10/sub_707/carry[1] ) );
  OA22X1 U6372 ( .IN1(n12696), .IN2(n13515), .IN3(n11444), .IN4(n11445), .Q(
        n11403) );
  NOR2X0 U6373 ( .IN1(n12697), .IN2(n13627), .QN(n11444) );
  NOR2X0 U6374 ( .IN1(\fadd_0_0_0_0_0/exponentdifferencexy [5]), .IN2(n12698), 
        .QN(n11446) );
  NOR2X0 U6375 ( .IN1(\fadd_0_0_0_0_4/exponentdifferencexy [5]), .IN2(n12738), 
        .QN(n11065) );
  NOR2X0 U6376 ( .IN1(\fadd_0_0_0_0_5/exponentdifferencexy [5]), .IN2(n12745), 
        .QN(n10984) );
  NOR2X0 U6377 ( .IN1(\fadd_0_0_0_0_2/exponentdifferencexy [5]), .IN2(n12718), 
        .QN(n11227) );
  NOR2X0 U6378 ( .IN1(\fadd_0_0_0_0_1/exponentdifferencexy [5]), .IN2(n12705), 
        .QN(n11363) );
  OA22X1 U6379 ( .IN1(n12736), .IN2(n13514), .IN3(n11063), .IN4(n11064), .Q(
        n11024) );
  NOR2X0 U6380 ( .IN1(n12737), .IN2(n13621), .QN(n11063) );
  OA22X1 U6381 ( .IN1(n12746), .IN2(n13511), .IN3(n10982), .IN4(n10983), .Q(
        n10943) );
  NOR2X0 U6382 ( .IN1(n12744), .IN2(n13624), .QN(n10982) );
  OA22X1 U6383 ( .IN1(n12716), .IN2(n13507), .IN3(n11225), .IN4(n11226), .Q(
        n11186) );
  NOR2X0 U6384 ( .IN1(n12717), .IN2(n13470), .QN(n11225) );
  OA22X1 U6385 ( .IN1(n12706), .IN2(n13509), .IN3(n11361), .IN4(n11362), .Q(
        n11322) );
  NOR2X0 U6386 ( .IN1(n12704), .IN2(n13622), .QN(n11361) );
  OA22X1 U6387 ( .IN1(n12776), .IN2(n13630), .IN3(n10739), .IN4(n10740), .Q(
        n10698) );
  NOR2X0 U6388 ( .IN1(n12774), .IN2(n13501), .QN(n10739) );
  NOR2X0 U6389 ( .IN1(\fadd_0_0_0_0_8/exponentdifferencexy [5]), .IN2(n12775), 
        .QN(n10741) );
  NOR2X0 U6390 ( .IN1(\fadd_0_0_0_0_9/exponentdifferencexy [5]), .IN2(n12785), 
        .QN(n10658) );
  NOR2X0 U6391 ( .IN1(\fadd_0_0_0_0_6/exponentdifferencexy [5]), .IN2(n12758), 
        .QN(n10903) );
  NOR2X0 U6392 ( .IN1(\fadd_0_0_0_0_7/exponentdifferencexy [5]), .IN2(n12765), 
        .QN(n10822) );
  NOR2X0 U6393 ( .IN1(\fadd_0_0_0_0_3/exponentdifferencexy [5]), .IN2(n12725), 
        .QN(n11146) );
  OA22X1 U6394 ( .IN1(n12786), .IN2(n13513), .IN3(n10656), .IN4(n10657), .Q(
        n10617) );
  NOR2X0 U6395 ( .IN1(n12784), .IN2(n13626), .QN(n10656) );
  OA22X1 U6396 ( .IN1(n12756), .IN2(n13508), .IN3(n10901), .IN4(n10902), .Q(
        n10862) );
  NOR2X0 U6397 ( .IN1(n12757), .IN2(n13471), .QN(n10901) );
  OA22X1 U6398 ( .IN1(n12766), .IN2(n13512), .IN3(n10820), .IN4(n10821), .Q(
        n10781) );
  NOR2X0 U6399 ( .IN1(n12764), .IN2(n13625), .QN(n10820) );
  OA22X1 U6400 ( .IN1(n12726), .IN2(n13510), .IN3(n11144), .IN4(n11145), .Q(
        n11105) );
  NOR2X0 U6401 ( .IN1(n12724), .IN2(n13623), .QN(n11144) );
  NOR2X0 U6402 ( .IN1(n12041), .IN2(n8850), .QN(n8839) );
  INVX0 U6403 ( .INP(n8787), .ZN(n14985) );
  NOR2X0 U6404 ( .IN1(n12067), .IN2(n14987), .QN(n8784) );
  NOR2X0 U6405 ( .IN1(n12028), .IN2(n12032), .QN(n11267) );
  NOR2X0 U6406 ( .IN1(n12032), .IN2(n8818), .QN(n8811) );
  NOR2X0 U6407 ( .IN1(n8850), .IN2(n13527), .QN(n8849) );
  NOR2X0 U6408 ( .IN1(n10558), .IN2(n12825), .QN(n10531) );
  NOR2X0 U6409 ( .IN1(n10531), .IN2(n10565), .QN(n10562) );
  NAND2X1 U6410 ( .IN1(n12068), .IN2(n14993), .QN(n8803) );
  NOR2X0 U6411 ( .IN1(n12821), .IN2(n12825), .QN(n10553) );
  NAND2X1 U6412 ( .IN1(n11609), .IN2(n14440), .QN(n13443) );
  NAND2X1 U6413 ( .IN1(n8842), .IN2(n8846), .QN(n8853) );
  OAI22X1 U6414 ( .IN1(n10698), .IN2(n11857), .IN3(n14311), .IN4(n11869), .QN(
        \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/n297_o[2] ) );
  NOR4X0 U6415 ( .IN1(n12001), .IN2(n12014), .IN3(n12015), .IN4(n12016), .QN(
        n8685) );
  OR3X1 U6416 ( .IN1(n15002), .IN2(n10675), .IN3(n14140), .Q(n10669) );
  AO221X1 U6417 ( .IN1(n14872), .IN2(\fadd_0_0_0_0_8/fracresultfar0 [0]), 
        .IN3(n10673), .IN4(\fadd_0_0_0_0_8/fracresultfar0 [1]), .IN5(n10674), 
        .Q(n14140) );
  NAND2X1 U6418 ( .IN1(n10663), .IN2(n10664), .QN(\fadd_0_0_0_0_8/round ) );
  NOR4X0 U6419 ( .IN1(n12169), .IN2(n12176), .IN3(n12177), .IN4(n12178), .QN(
        n9070) );
  OR3X1 U6420 ( .IN1(n14956), .IN2(n11001), .IN3(n14141), .Q(n10995) );
  AO221X1 U6421 ( .IN1(n14777), .IN2(\fadd_0_0_0_0_4/fracresultfar0 [0]), 
        .IN3(n10999), .IN4(\fadd_0_0_0_0_4/fracresultfar0 [1]), .IN5(n11000), 
        .Q(n14141) );
  NAND2X1 U6422 ( .IN1(n10989), .IN2(n10990), .QN(\fadd_0_0_0_0_4/round ) );
  NOR4X0 U6423 ( .IN1(n12291), .IN2(n12297), .IN3(n12298), .IN4(n12299), .QN(
        n9290) );
  OR3X1 U6424 ( .IN1(n14946), .IN2(n11163), .IN3(n14142), .Q(n11157) );
  AO221X1 U6425 ( .IN1(n14724), .IN2(\fadd_0_0_0_0_2/fracresultfar0 [0]), 
        .IN3(n11161), .IN4(\fadd_0_0_0_0_2/fracresultfar0 [1]), .IN5(n11162), 
        .Q(n14142) );
  NAND2X1 U6426 ( .IN1(n11151), .IN2(n11152), .QN(\fadd_0_0_0_0_2/round ) );
  INVX0 U6427 ( .INP(n8678), .ZN(n14859) );
  INVX0 U6428 ( .INP(n9065), .ZN(n14764) );
  INVX0 U6429 ( .INP(n9285), .ZN(n14711) );
  NOR2X0 U6430 ( .IN1(n12825), .IN2(n12820), .QN(n10559) );
  NOR2X0 U6431 ( .IN1(n12824), .IN2(n10538), .QN(n10536) );
  OAI22X1 U6432 ( .IN1(n14917), .IN2(n11999), .IN3(n14860), .IN4(n12827), .QN(
        n12412) );
  NOR2X0 U6433 ( .IN1(n12820), .IN2(n12824), .QN(n10538) );
  OAI22X1 U6434 ( .IN1(n14184), .IN2(n12004), .IN3(n8245), .IN4(n12827), .QN(
        n12417) );
  NOR2X0 U6435 ( .IN1(n12821), .IN2(n12824), .QN(n10550) );
  NOR2X0 U6436 ( .IN1(n11924), .IN2(n12824), .QN(n10540) );
  NOR2X0 U6437 ( .IN1(n12821), .IN2(n12823), .QN(n10564) );
  NOR4X0 U6438 ( .IN1(n12203), .IN2(n12207), .IN3(n12208), .IN4(n12209), .QN(
        n9141) );
  INVX0 U6439 ( .INP(\fadd_0_0_0_0_6/resultrounded [9]), .ZN(n14816) );
  NOR4X0 U6440 ( .IN1(n12140), .IN2(n12146), .IN3(n12147), .IN4(n12148), .QN(
        n8960) );
  INVX0 U6441 ( .INP(\fadd_0_0_0_0_0/resultrounded [9]), .ZN(n14668) );
  OR3X1 U6442 ( .IN1(n14958), .IN2(n11380), .IN3(n14143), .Q(n11374) );
  AO221X1 U6443 ( .IN1(n14671), .IN2(\fadd_0_0_0_0_0/fracresultfar0 [0]), 
        .IN3(n11378), .IN4(\fadd_0_0_0_0_0/fracresultfar0 [1]), .IN5(n11379), 
        .Q(n14143) );
  OR3X1 U6444 ( .IN1(n14953), .IN2(n10839), .IN3(n14144), .Q(n10833) );
  AO221X1 U6445 ( .IN1(n14819), .IN2(\fadd_0_0_0_0_6/fracresultfar0 [0]), 
        .IN3(n10837), .IN4(\fadd_0_0_0_0_6/fracresultfar0 [1]), .IN5(n10838), 
        .Q(n14144) );
  NAND2X1 U6446 ( .IN1(n11368), .IN2(n11369), .QN(\fadd_0_0_0_0_0/round ) );
  NAND2X1 U6447 ( .IN1(n10827), .IN2(n10828), .QN(\fadd_0_0_0_0_6/round ) );
  NOR4X0 U6448 ( .IN1(n12231), .IN2(n12237), .IN3(n12238), .IN4(n12239), .QN(
        n9204) );
  INVX0 U6449 ( .INP(\fadd_0_0_0_0_7/resultrounded [9]), .ZN(n14837) );
  NOR4X0 U6450 ( .IN1(n12261), .IN2(n12267), .IN3(n12268), .IN4(n12269), .QN(
        n9246) );
  INVX0 U6451 ( .INP(\fadd_0_0_0_0_5/resultrounded [9]), .ZN(n14795) );
  OR3X1 U6452 ( .IN1(n14951), .IN2(n10758), .IN3(n14145), .Q(n10752) );
  AO221X1 U6453 ( .IN1(n14840), .IN2(\fadd_0_0_0_0_7/fracresultfar0 [0]), 
        .IN3(n10756), .IN4(\fadd_0_0_0_0_7/fracresultfar0 [1]), .IN5(n10757), 
        .Q(n14145) );
  OR3X1 U6454 ( .IN1(n14949), .IN2(n10920), .IN3(n14146), .Q(n10914) );
  AO221X1 U6455 ( .IN1(n14798), .IN2(\fadd_0_0_0_0_5/fracresultfar0 [0]), 
        .IN3(n10918), .IN4(\fadd_0_0_0_0_5/fracresultfar0 [1]), .IN5(n10919), 
        .Q(n14146) );
  NAND2X1 U6456 ( .IN1(n10746), .IN2(n10747), .QN(\fadd_0_0_0_0_7/round ) );
  NAND2X1 U6457 ( .IN1(n10908), .IN2(n10909), .QN(\fadd_0_0_0_0_5/round ) );
  OR3X1 U6458 ( .IN1(n14960), .IN2(n10594), .IN3(n14147), .Q(n10588) );
  AO221X1 U6459 ( .IN1(n14893), .IN2(\fadd_0_0_0_0_9/fracresultfar0 [0]), 
        .IN3(n10592), .IN4(\fadd_0_0_0_0_9/fracresultfar0 [1]), .IN5(n10593), 
        .Q(n14147) );
  OR3X1 U6460 ( .IN1(n14947), .IN2(n11082), .IN3(n14148), .Q(n11076) );
  AO221X1 U6461 ( .IN1(n14745), .IN2(\fadd_0_0_0_0_3/fracresultfar0 [0]), 
        .IN3(n11080), .IN4(\fadd_0_0_0_0_3/fracresultfar0 [1]), .IN5(n11081), 
        .Q(n14148) );
  OR3X1 U6462 ( .IN1(n14942), .IN2(n11299), .IN3(n14149), .Q(n11293) );
  AO221X1 U6463 ( .IN1(n14692), .IN2(\fadd_0_0_0_0_1/fracresultfar0 [0]), 
        .IN3(n11297), .IN4(\fadd_0_0_0_0_1/fracresultfar0 [1]), .IN5(n11298), 
        .Q(n14149) );
  NOR4X0 U6464 ( .IN1(n12095), .IN2(n12102), .IN3(n12103), .IN4(n12104), .QN(
        n8912) );
  INVX0 U6465 ( .INP(\fadd_0_0_0_0_9/resultrounded [9]), .ZN(n14890) );
  NOR4X0 U6466 ( .IN1(n12320), .IN2(n12327), .IN3(n12328), .IN4(n12329), .QN(
        n9352) );
  INVX0 U6467 ( .INP(\fadd_0_0_0_0_3/resultrounded [9]), .ZN(n14742) );
  NOR4X0 U6468 ( .IN1(n12351), .IN2(n12359), .IN3(n12360), .IN4(n12361), .QN(
        n9394) );
  INVX0 U6469 ( .INP(\fadd_0_0_0_0_1/resultrounded [9]), .ZN(n14689) );
  NAND2X1 U6470 ( .IN1(n10582), .IN2(n10583), .QN(\fadd_0_0_0_0_9/round ) );
  NAND2X1 U6471 ( .IN1(n11070), .IN2(n11071), .QN(\fadd_0_0_0_0_3/round ) );
  NAND2X1 U6472 ( .IN1(n11287), .IN2(n11288), .QN(\fadd_0_0_0_0_1/round ) );
  NOR2X0 U6473 ( .IN1(n12822), .IN2(n12823), .QN(n10555) );
  OAI22X1 U6474 ( .IN1(n14917), .IN2(n11971), .IN3(n14861), .IN4(n12827), .QN(
        n12377) );
  XOR2X1 U6475 ( .IN1(n14182), .IN2(n14150), .Q(
        \fmul_0_0_0_0_10/roundingadder/add_1_root_add_57/SUM[10] ) );
  NAND2X1 U6476 ( .IN1(n14158), .IN2(
        \fmul_0_0_0_0_10/roundingadder/add_1_root_add_57/A[9] ), .QN(n14182)
         );
  AND2X1 U6477 ( .IN1(\fmul_0_0_0_0_10/roundingadder/add_1_root_add_57/A[0] ), 
        .IN2(\fmul_0_0_0_0_10/roundingadder/add_1_root_add_57/CI ), .Q(n14151)
         );
  AND2X1 U6478 ( .IN1(\fmul_0_0_0_0_10/roundingadder/add_1_root_add_57/A[1] ), 
        .IN2(n14151), .Q(n14152) );
  AND2X1 U6479 ( .IN1(\fmul_0_0_0_0_10/roundingadder/add_1_root_add_57/A[2] ), 
        .IN2(n14152), .Q(n14153) );
  AND2X1 U6480 ( .IN1(\fmul_0_0_0_0_10/roundingadder/add_1_root_add_57/A[3] ), 
        .IN2(n14153), .Q(n14154) );
  AND2X1 U6481 ( .IN1(\fmul_0_0_0_0_10/roundingadder/add_1_root_add_57/A[4] ), 
        .IN2(n14154), .Q(n14155) );
  AND2X1 U6482 ( .IN1(\fmul_0_0_0_0_10/roundingadder/add_1_root_add_57/A[5] ), 
        .IN2(n14155), .Q(n14156) );
  AND2X1 U6483 ( .IN1(\fmul_0_0_0_0_10/roundingadder/add_1_root_add_57/A[7] ), 
        .IN2(n14160), .Q(n14157) );
  AND2X1 U6484 ( .IN1(\fmul_0_0_0_0_10/roundingadder/add_1_root_add_57/A[8] ), 
        .IN2(n14157), .Q(n14158) );
  OR2X1 U6485 ( .IN1(n11958), .IN2(n14159), .Q(n8887) );
  AND3X1 U6486 ( .IN1(n14961), .IN2(n13771), .IN3(
        \fmul_0_0_0_0_10/roundingadder/add_1_root_add_57/SUM[9] ), .Q(n14159)
         );
  AND2X1 U6487 ( .IN1(\fmul_0_0_0_0_10/roundingadder/add_1_root_add_57/A[6] ), 
        .IN2(n14156), .Q(n14160) );
  NOR2X0 U6488 ( .IN1(n11924), .IN2(n13499), .QN(n10542) );
  INVX0 U6489 ( .INP(n10519), .ZN(n14924) );
  NAND2X1 U6490 ( .IN1(n12820), .IN2(n12824), .QN(n10544) );
  OAI22X1 U6491 ( .IN1(n14184), .IN2(n11975), .IN3(n14862), .IN4(n12827), .QN(
        n12382) );
  NOR2X0 U6492 ( .IN1(\fmul_0_0_0_0_10/roundingadder/add_1_root_add_57/SUM[9] ), .IN2(\fmul_0_0_0_0_10/roundingadder/add_1_root_add_57/SUM[10] ), .QN(n8894)
         );
  OAI22X1 U6493 ( .IN1(n10698), .IN2(n11859), .IN3(n14311), .IN4(n11871), .QN(
        \fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/n297_o[4] ) );
  OAI22X1 U6494 ( .IN1(n14184), .IN2(n11979), .IN3(n14863), .IN4(n12827), .QN(
        n12387) );
  OAI22X1 U6495 ( .IN1(n14917), .IN2(n11983), .IN3(n14864), .IN4(n12827), .QN(
        n12392) );
  OAI22X1 U6496 ( .IN1(n14184), .IN2(n11987), .IN3(n14865), .IN4(n12827), .QN(
        n12397) );
  INVX0 U6497 ( .INP(n10400), .ZN(n14913) );
  NAND2X1 U6498 ( .IN1(n11927), .IN2(n12832), .QN(n10400) );
  OR2X1 U6499 ( .IN1(n14161), .IN2(n10402), .Q(n10397) );
  OAI22X1 U6500 ( .IN1(n14917), .IN2(n11991), .IN3(n14866), .IN4(n12827), .QN(
        n12402) );
  NAND2X1 U6501 ( .IN1(n11924), .IN2(n12823), .QN(n10518) );
  OAI22X1 U6502 ( .IN1(n14184), .IN2(n11995), .IN3(n14867), .IN4(n12827), .QN(
        n12407) );
  OAI22X1 U6503 ( .IN1(n14184), .IN2(n11967), .IN3(n14868), .IN4(n12827), .QN(
        n12372) );
  OAI22X1 U6504 ( .IN1(n14917), .IN2(n11963), .IN3(n14869), .IN4(n12827), .QN(
        n12367) );
  OR3X1 U6505 ( .IN1(n14162), .IN2(n14163), .IN3(n8988), .Q(n8947) );
  AND2X1 U6506 ( .IN1(n8989), .IN2(n8990), .Q(n14163) );
  NOR2X0 U6507 ( .IN1(n12068), .IN2(n12061), .QN(n8856) );
  NOR2X0 U6508 ( .IN1(\fmul_0_0_0_0_0/expsigpostround [9]), .IN2(
        \fmul_0_0_0_0_0/expsigpostround [10]), .QN(n9003) );
  NAND2X1 U6509 ( .IN1(n12822), .IN2(n12820), .QN(n10493) );
  NOR2X0 U6510 ( .IN1(n10485), .IN2(n10486), .QN(\fmul_0_0_0_0_10/n98 ) );
  NOR2X0 U6511 ( .IN1(n12822), .IN2(n12825), .QN(n10491) );
  NOR2X0 U6512 ( .IN1(\fadd_0_0_0_0_8/exponentdifferenceyx [3]), .IN2(
        \fadd_0_0_0_0_8/exponentdifferenceyx [4]), .QN(n10701) );
  XOR3X1 U6513 ( .IN1(n5410), .IN2(n14624), .IN3(
        \fadd_0_0_0_0_8/sub_710/carry [4]), .Q(
        \fadd_0_0_0_0_8/exponentdifferenceyx [4]) );
  NOR2X0 U6514 ( .IN1(\fadd_0_0_0_0_9/exponentdifferenceyx [3]), .IN2(
        \fadd_0_0_0_0_9/exponentdifferenceyx [4]), .QN(n10620) );
  XOR3X1 U6515 ( .IN1(n5338), .IN2(n14635), .IN3(
        \fadd_0_0_0_0_9/sub_710/carry [4]), .Q(
        \fadd_0_0_0_0_9/exponentdifferenceyx [4]) );
  NOR2X0 U6516 ( .IN1(\fadd_0_0_0_0_7/exponentdifferenceyx [3]), .IN2(
        \fadd_0_0_0_0_7/exponentdifferenceyx [4]), .QN(n10784) );
  XOR3X1 U6517 ( .IN1(n5482), .IN2(n14613), .IN3(
        \fadd_0_0_0_0_7/sub_710/carry [4]), .Q(
        \fadd_0_0_0_0_7/exponentdifferenceyx [4]) );
  NOR2X0 U6518 ( .IN1(\fadd_0_0_0_0_0/exponentdifferenceyx [3]), .IN2(
        \fadd_0_0_0_0_0/exponentdifferenceyx [4]), .QN(n11406) );
  XOR3X1 U6519 ( .IN1(n5986), .IN2(n14536), .IN3(
        \fadd_0_0_0_0_0/sub_710/carry [4]), .Q(
        \fadd_0_0_0_0_0/exponentdifferenceyx [4]) );
  NOR2X0 U6520 ( .IN1(\fadd_0_0_0_0_4/exponentdifferenceyx [3]), .IN2(
        \fadd_0_0_0_0_4/exponentdifferenceyx [4]), .QN(n11027) );
  XOR3X1 U6521 ( .IN1(n5698), .IN2(n14580), .IN3(
        \fadd_0_0_0_0_4/sub_710/carry [4]), .Q(
        \fadd_0_0_0_0_4/exponentdifferenceyx [4]) );
  NOR2X0 U6522 ( .IN1(\fadd_0_0_0_0_6/exponentdifferenceyx [3]), .IN2(
        \fadd_0_0_0_0_6/exponentdifferenceyx [4]), .QN(n10865) );
  XOR3X1 U6523 ( .IN1(n5554), .IN2(n14602), .IN3(
        \fadd_0_0_0_0_6/sub_710/carry [4]), .Q(
        \fadd_0_0_0_0_6/exponentdifferenceyx [4]) );
  NOR2X0 U6524 ( .IN1(\fadd_0_0_0_0_5/exponentdifferenceyx [3]), .IN2(
        \fadd_0_0_0_0_5/exponentdifferenceyx [4]), .QN(n10946) );
  XOR3X1 U6525 ( .IN1(n5626), .IN2(n14591), .IN3(
        \fadd_0_0_0_0_5/sub_710/carry [4]), .Q(
        \fadd_0_0_0_0_5/exponentdifferenceyx [4]) );
  NOR2X0 U6526 ( .IN1(\fadd_0_0_0_0_3/exponentdifferenceyx [3]), .IN2(
        \fadd_0_0_0_0_3/exponentdifferenceyx [4]), .QN(n11108) );
  XOR3X1 U6527 ( .IN1(n5770), .IN2(n14569), .IN3(
        \fadd_0_0_0_0_3/sub_710/carry [4]), .Q(
        \fadd_0_0_0_0_3/exponentdifferenceyx [4]) );
  NOR2X0 U6528 ( .IN1(\fadd_0_0_0_0_2/exponentdifferenceyx [3]), .IN2(
        \fadd_0_0_0_0_2/exponentdifferenceyx [4]), .QN(n11189) );
  XOR3X1 U6529 ( .IN1(n5842), .IN2(n14562), .IN3(
        \fadd_0_0_0_0_2/sub_710/carry [4]), .Q(
        \fadd_0_0_0_0_2/exponentdifferenceyx [4]) );
  NOR2X0 U6530 ( .IN1(\fadd_0_0_0_0_1/exponentdifferenceyx [3]), .IN2(
        \fadd_0_0_0_0_1/exponentdifferenceyx [4]), .QN(n11325) );
  XOR3X1 U6531 ( .IN1(n5914), .IN2(n14547), .IN3(
        \fadd_0_0_0_0_1/sub_710/carry [4]), .Q(
        \fadd_0_0_0_0_1/exponentdifferenceyx [4]) );
  NOR2X0 U6532 ( .IN1(n14186), .IN2(n12832), .QN(n9451) );
  NAND2X1 U6533 ( .IN1(n13635), .IN2(n14179), .QN(
        \fadd_0_0_0_0_10/sub_710/carry[1] ) );
  NOR2X0 U6534 ( .IN1(n10397), .IN2(n12836), .QN(n9446) );
  NOR2X0 U6535 ( .IN1(n12865), .IN2(n12846), .QN(n10680) );
  NOR2X0 U6536 ( .IN1(n12857), .IN2(n12842), .QN(n11006) );
  NOR2X0 U6537 ( .IN1(n12853), .IN2(n12840), .QN(n11168) );
  NAND2X1 U6538 ( .IN1(n14178), .IN2(n13714), .QN(
        \fadd_0_0_0_0_10/sub_784/carry[1] ) );
  INVX0 U6539 ( .INP(\fadd_0_0_0_0_10/norm/U5/Z_5 ), .ZN(n14178) );
  NOR2X0 U6540 ( .IN1(\fmul_0_0_0_0_1/expsigpostround [9]), .IN2(
        \fmul_0_0_0_0_1/expsigpostround [10]), .QN(n9419) );
  NOR2X0 U6541 ( .IN1(\fmul_0_0_0_0_9/expsigpostround [9]), .IN2(
        \fmul_0_0_0_0_9/expsigpostround [10]), .QN(n8936) );
  NOR2X0 U6542 ( .IN1(\fmul_0_0_0_0_7/expsigpostround [9]), .IN2(
        \fmul_0_0_0_0_7/expsigpostround [10]), .QN(n9228) );
  NOR2X0 U6543 ( .IN1(\fmul_0_0_0_0_5/expsigpostround [9]), .IN2(
        \fmul_0_0_0_0_5/expsigpostround [10]), .QN(n9270) );
  NOR2X0 U6544 ( .IN1(\fmul_0_0_0_0_3/expsigpostround [9]), .IN2(
        \fmul_0_0_0_0_3/expsigpostround [10]), .QN(n9376) );
  OR2X1 U6545 ( .IN1(n11941), .IN2(n14164), .Q(n9369) );
  AND3X1 U6546 ( .IN1(n14897), .IN2(n13767), .IN3(
        \fmul_0_0_0_0_3/expsigpostround [9]), .Q(n14164) );
  OR2X1 U6547 ( .IN1(n11956), .IN2(n14165), .Q(n8929) );
  AND3X1 U6548 ( .IN1(n14903), .IN2(n13770), .IN3(
        \fmul_0_0_0_0_9/expsigpostround [9]), .Q(n14165) );
  OR2X1 U6549 ( .IN1(n11947), .IN2(n14166), .Q(n9221) );
  AND3X1 U6550 ( .IN1(n14901), .IN2(n13769), .IN3(
        \fmul_0_0_0_0_7/expsigpostround [9]), .Q(n14166) );
  OR2X1 U6551 ( .IN1(n11945), .IN2(n14167), .Q(n9263) );
  AND3X1 U6552 ( .IN1(n14899), .IN2(n13768), .IN3(
        \fmul_0_0_0_0_5/expsigpostround [9]), .Q(n14167) );
  OR2X1 U6553 ( .IN1(n11939), .IN2(n14168), .Q(n9412) );
  AND3X1 U6554 ( .IN1(n14895), .IN2(n13766), .IN3(
        \fmul_0_0_0_0_1/expsigpostround [9]), .Q(n14168) );
  NOR2X0 U6555 ( .IN1(n11921), .IN2(n14937), .QN(n8669) );
  NOR2X0 U6556 ( .IN1(n11917), .IN2(n14936), .QN(n8665) );
  NOR2X0 U6557 ( .IN1(n11913), .IN2(n14935), .QN(n8661) );
  NOR2X0 U6558 ( .IN1(n11909), .IN2(n14934), .QN(n8657) );
  NOR2X0 U6559 ( .IN1(n11905), .IN2(n14933), .QN(n8653) );
  NOR2X0 U6560 ( .IN1(n11901), .IN2(n14932), .QN(n8649) );
  NOR2X0 U6561 ( .IN1(n11897), .IN2(n14931), .QN(n8645) );
  NOR2X0 U6562 ( .IN1(n11893), .IN2(n14930), .QN(n8641) );
  NOR2X0 U6563 ( .IN1(n11885), .IN2(n14929), .QN(n8637) );
  NOR2X0 U6564 ( .IN1(n11881), .IN2(n14928), .QN(n8633) );
  NOR2X0 U6565 ( .IN1(n10419), .IN2(n11598), .QN(n8668) );
  NOR2X0 U6566 ( .IN1(n10418), .IN2(n11585), .QN(n8664) );
  NOR2X0 U6567 ( .IN1(n10417), .IN2(n11572), .QN(n8660) );
  NOR2X0 U6568 ( .IN1(n10416), .IN2(n11559), .QN(n8656) );
  NOR2X0 U6569 ( .IN1(n10415), .IN2(n11546), .QN(n8652) );
  NOR2X0 U6570 ( .IN1(n10414), .IN2(n11533), .QN(n8648) );
  NOR2X0 U6571 ( .IN1(n10413), .IN2(n11520), .QN(n8644) );
  NOR2X0 U6572 ( .IN1(n10412), .IN2(n11507), .QN(n8640) );
  NOR2X0 U6573 ( .IN1(n10411), .IN2(n11485), .QN(n8636) );
  NOR2X0 U6574 ( .IN1(n10410), .IN2(n11472), .QN(n8632) );
  NOR2X0 U6575 ( .IN1(n10402), .IN2(n12835), .QN(n9452) );
  NAND2X1 U6576 ( .IN1(n12830), .IN2(n11928), .QN(n10393) );
  NOR2X0 U6577 ( .IN1(n12849), .IN2(n12838), .QN(n11385) );
  NOR2X0 U6578 ( .IN1(n12861), .IN2(n12844), .QN(n10844) );
  NOR2X0 U6579 ( .IN1(n12863), .IN2(n12845), .QN(n10763) );
  NOR2X0 U6580 ( .IN1(n12859), .IN2(n12843), .QN(n10925) );
  NOR2X0 U6581 ( .IN1(n12867), .IN2(n12847), .QN(n10599) );
  NOR2X0 U6582 ( .IN1(n12855), .IN2(n12841), .QN(n11087) );
  NOR2X0 U6583 ( .IN1(n12851), .IN2(n12839), .QN(n11304) );
  NOR2X0 U6584 ( .IN1(n10400), .IN2(n12833), .QN(n9454) );
  NOR2X0 U6585 ( .IN1(n10393), .IN2(n12831), .QN(n9443) );
  NOR2X0 U6586 ( .IN1(n13497), .IN2(n12826), .QN(n8732) );
  INVX0 U6587 ( .INP(\fmul_0_0_0_0_0/expsigpostround [10]), .ZN(n14894) );
  INVX0 U6588 ( .INP(\fmul_0_0_0_0_8/expsigpostround[10] ), .ZN(n14902) );
  XOR2X1 U6589 ( .IN1(
        \add_1_root_fmul_0_0_0_0_8/roundingadder/add_57/carry [9]), .IN2(
        n14170), .Q(n14169) );
  NOR2X0 U6590 ( .IN1(n11598), .IN2(n10626), .QN(
        \fadd_0_0_0_0_9/norm/level1 [1]) );
  NOR2X0 U6591 ( .IN1(n11585), .IN2(n10707), .QN(
        \fadd_0_0_0_0_8/norm/level1 [1]) );
  NOR2X0 U6592 ( .IN1(n11572), .IN2(n10790), .QN(
        \fadd_0_0_0_0_7/norm/level1 [1]) );
  NOR2X0 U6593 ( .IN1(n11559), .IN2(n10871), .QN(
        \fadd_0_0_0_0_6/norm/level1 [1]) );
  NOR2X0 U6594 ( .IN1(n11546), .IN2(n10952), .QN(
        \fadd_0_0_0_0_5/norm/level1 [1]) );
  NOR2X0 U6595 ( .IN1(n11533), .IN2(n11033), .QN(
        \fadd_0_0_0_0_4/norm/level1 [1]) );
  NOR2X0 U6596 ( .IN1(n11520), .IN2(n11114), .QN(
        \fadd_0_0_0_0_3/norm/level1 [1]) );
  NOR2X0 U6597 ( .IN1(n11507), .IN2(n11195), .QN(
        \fadd_0_0_0_0_2/norm/level1 [1]) );
  NOR2X0 U6598 ( .IN1(n11485), .IN2(n11331), .QN(
        \fadd_0_0_0_0_1/norm/level1 [1]) );
  NOR2X0 U6599 ( .IN1(n11472), .IN2(n11412), .QN(
        \fadd_0_0_0_0_0/norm/level1 [1]) );
  NOR2X0 U6600 ( .IN1(n11597), .IN2(n10626), .QN(
        \fadd_0_0_0_0_9/norm/level1 [0]) );
  NOR2X0 U6601 ( .IN1(n11584), .IN2(n10707), .QN(
        \fadd_0_0_0_0_8/norm/level1 [0]) );
  NOR2X0 U6602 ( .IN1(n11571), .IN2(n10790), .QN(
        \fadd_0_0_0_0_7/norm/level1 [0]) );
  NOR2X0 U6603 ( .IN1(n11558), .IN2(n10871), .QN(
        \fadd_0_0_0_0_6/norm/level1 [0]) );
  NOR2X0 U6604 ( .IN1(n11545), .IN2(n10952), .QN(
        \fadd_0_0_0_0_5/norm/level1 [0]) );
  NOR2X0 U6605 ( .IN1(n11532), .IN2(n11033), .QN(
        \fadd_0_0_0_0_4/norm/level1 [0]) );
  NOR2X0 U6606 ( .IN1(n11519), .IN2(n11114), .QN(
        \fadd_0_0_0_0_3/norm/level1 [0]) );
  NOR2X0 U6607 ( .IN1(n11506), .IN2(n11195), .QN(
        \fadd_0_0_0_0_2/norm/level1 [0]) );
  NOR2X0 U6608 ( .IN1(n11484), .IN2(n11331), .QN(
        \fadd_0_0_0_0_1/norm/level1 [0]) );
  NOR2X0 U6609 ( .IN1(n11471), .IN2(n11412), .QN(
        \fadd_0_0_0_0_0/norm/level1 [0]) );
  NAND4X0 U6610 ( .IN1(n12014), .IN2(n12015), .IN3(n12016), .IN4(n13723), .QN(
        n8683) );
  NAND4X0 U6611 ( .IN1(n12176), .IN2(n12177), .IN3(n12178), .IN4(n13725), .QN(
        n9068) );
  NAND4X0 U6612 ( .IN1(n12297), .IN2(n12298), .IN3(n12299), .IN4(n13727), .QN(
        n9288) );
  NAND2X1 U6613 ( .IN1(n11952), .IN2(n14917), .QN(n8999) );
  NAND2X1 U6614 ( .IN1(\fadd_0_0_0_0_8/syncx_d2 [9]), .IN2(n8690), .QN(n8689)
         );
  NOR2X0 U6615 ( .IN1(n12016), .IN2(n13735), .QN(n8691) );
  INVX0 U6616 ( .INP(n8247), .ZN(n15000) );
  NAND2X1 U6617 ( .IN1(\fadd_0_0_0_0_4/syncx_d2 [9]), .IN2(n9075), .QN(n9074)
         );
  NOR2X0 U6618 ( .IN1(n12178), .IN2(n13737), .QN(n9076) );
  NAND2X1 U6619 ( .IN1(\fadd_0_0_0_0_2/syncx_d2 [9]), .IN2(n9294), .QN(n9293)
         );
  NOR2X0 U6620 ( .IN1(n11498), .IN2(n11238), .QN(\fadd_0_0_0_0_10/norm/U5/Z_0 ) );
  NOR2X0 U6621 ( .IN1(n11499), .IN2(n11238), .QN(\fadd_0_0_0_0_10/norm/U5/Z_1 ) );
  NOR2X0 U6622 ( .IN1(n13727), .IN2(\fadd_0_0_0_0_2/syncsigny_d2 ), .QN(n9296)
         );
  OAI22X1 U6623 ( .IN1(n14184), .IN2(n12010), .IN3(n8247), .IN4(n12827), .QN(
        n12422) );
  NAND4X0 U6624 ( .IN1(n12102), .IN2(n12103), .IN3(n12104), .IN4(n13732), .QN(
        n8910) );
  NAND4X0 U6625 ( .IN1(n12327), .IN2(n12328), .IN3(n12329), .IN4(n13731), .QN(
        n9350) );
  NAND4X0 U6626 ( .IN1(n12359), .IN2(n12360), .IN3(n12361), .IN4(n13730), .QN(
        n9392) );
  NAND2X1 U6627 ( .IN1(\fadd_0_0_0_0_9/syncx_d2 [9]), .IN2(n8916), .QN(n8915)
         );
  NOR2X0 U6628 ( .IN1(n12104), .IN2(n13739), .QN(n8917) );
  NAND2X1 U6629 ( .IN1(\fadd_0_0_0_0_3/syncx_d2 [9]), .IN2(n9356), .QN(n9355)
         );
  NOR2X0 U6630 ( .IN1(n12329), .IN2(n13740), .QN(n9357) );
  NAND2X1 U6631 ( .IN1(\fadd_0_0_0_0_1/syncx_d2 [9]), .IN2(n9398), .QN(n9397)
         );
  NOR2X0 U6632 ( .IN1(n12361), .IN2(n13741), .QN(n9399) );
  NAND2X1 U6633 ( .IN1(\fadd_0_0_0_0_0/syncx_d2 [9]), .IN2(n8965), .QN(n8964)
         );
  NAND2X1 U6634 ( .IN1(\fadd_0_0_0_0_7/syncx_d2 [9]), .IN2(n9208), .QN(n9207)
         );
  NAND2X1 U6635 ( .IN1(\fadd_0_0_0_0_5/syncx_d2 [9]), .IN2(n9250), .QN(n9249)
         );
  NAND2X1 U6636 ( .IN1(\fadd_0_0_0_0_6/syncx_d2 [9]), .IN2(n9145), .QN(n9144)
         );
  NAND2X1 U6637 ( .IN1(\fadd_0_0_0_0_10/U12/DATA3_0 ), .IN2(n8794), .QN(n8793)
         );
  NOR2X0 U6638 ( .IN1(n13729), .IN2(\fadd_0_0_0_0_0/syncsigny_d2 ), .QN(n8967)
         );
  NOR2X0 U6639 ( .IN1(n13724), .IN2(\fadd_0_0_0_0_10/n147 ), .QN(n8796) );
  NOR2X0 U6640 ( .IN1(n13734), .IN2(\fadd_0_0_0_0_7/syncsigny_d2 ), .QN(n9210)
         );
  NOR2X0 U6641 ( .IN1(n13733), .IN2(\fadd_0_0_0_0_5/syncsigny_d2 ), .QN(n9252)
         );
  NOR2X0 U6642 ( .IN1(n13728), .IN2(\fadd_0_0_0_0_6/syncsigny_d2 ), .QN(n9147)
         );
  NAND2X1 U6643 ( .IN1(n11655), .IN2(n12815), .QN(\fmul_0_0_0_0_10/U9/Z_1 ) );
  NAND2X1 U6644 ( .IN1(n11651), .IN2(n12787), .QN(\fmul_0_0_0_0_9/exc [1]) );
  NAND2X1 U6645 ( .IN1(n11647), .IN2(n12777), .QN(\fmul_0_0_0_0_8/exc [1]) );
  NAND2X1 U6646 ( .IN1(n11643), .IN2(n12767), .QN(\fmul_0_0_0_0_7/exc [1]) );
  NAND2X1 U6647 ( .IN1(n11639), .IN2(n12749), .QN(\fmul_0_0_0_0_6/exc [1]) );
  NAND2X1 U6648 ( .IN1(n11635), .IN2(n12747), .QN(\fmul_0_0_0_0_5/exc [1]) );
  NAND2X1 U6649 ( .IN1(n11631), .IN2(n12729), .QN(\fmul_0_0_0_0_4/exc [1]) );
  NAND2X1 U6650 ( .IN1(n11627), .IN2(n12727), .QN(\fmul_0_0_0_0_3/exc [1]) );
  NAND2X1 U6651 ( .IN1(n11623), .IN2(n12709), .QN(\fmul_0_0_0_0_2/exc [1]) );
  NAND2X1 U6652 ( .IN1(n11619), .IN2(n12707), .QN(\fmul_0_0_0_0_1/exc [1]) );
  NAND2X1 U6653 ( .IN1(n11615), .IN2(n12689), .QN(\fmul_0_0_0_0_0/exc [1]) );
  NAND2X1 U6654 ( .IN1(n12697), .IN2(n12696), .QN(\fadd_0_0_0_0_0/newx [11])
         );
  NAND2X1 U6655 ( .IN1(n12802), .IN2(n12808), .QN(\fadd_0_0_0_0_10/U29/Z_11 )
         );
  NAND2X1 U6656 ( .IN1(n12774), .IN2(n12776), .QN(\fadd_0_0_0_0_8/newx [11])
         );
  NAND2X1 U6657 ( .IN1(n11589), .IN2(n11590), .QN(n10678) );
  NAND2X1 U6658 ( .IN1(n11591), .IN2(n11592), .QN(n10677) );
  NAND2X1 U6659 ( .IN1(n11500), .IN2(n11501), .QN(n11233) );
  NAND2X1 U6660 ( .IN1(n11502), .IN2(n11503), .QN(n11232) );
  NAND2X1 U6661 ( .IN1(n11602), .IN2(n11603), .QN(n10597) );
  NAND2X1 U6662 ( .IN1(n11604), .IN2(n11605), .QN(n10596) );
  NAND2X1 U6663 ( .IN1(n11476), .IN2(n11477), .QN(n11383) );
  NAND2X1 U6664 ( .IN1(n11478), .IN2(n11479), .QN(n11382) );
  NAND2X1 U6665 ( .IN1(n11537), .IN2(n11538), .QN(n11004) );
  NAND2X1 U6666 ( .IN1(n11539), .IN2(n11540), .QN(n11003) );
  NAND2X1 U6667 ( .IN1(n11563), .IN2(n11564), .QN(n10842) );
  NAND2X1 U6668 ( .IN1(n11565), .IN2(n11566), .QN(n10841) );
  NAND2X1 U6669 ( .IN1(n11576), .IN2(n11577), .QN(n10761) );
  NAND2X1 U6670 ( .IN1(n11578), .IN2(n11579), .QN(n10760) );
  NAND2X1 U6671 ( .IN1(n11550), .IN2(n11551), .QN(n10923) );
  NAND2X1 U6672 ( .IN1(n11552), .IN2(n11553), .QN(n10922) );
  NAND2X1 U6673 ( .IN1(n11524), .IN2(n11525), .QN(n11085) );
  NAND2X1 U6674 ( .IN1(n11526), .IN2(n11527), .QN(n11084) );
  NAND2X1 U6675 ( .IN1(n11511), .IN2(n11512), .QN(n11166) );
  NAND2X1 U6676 ( .IN1(n11513), .IN2(n11514), .QN(n11165) );
  NAND2X1 U6677 ( .IN1(n11489), .IN2(n11490), .QN(n11302) );
  NAND2X1 U6678 ( .IN1(n11491), .IN2(n11492), .QN(n11301) );
  NAND2X1 U6679 ( .IN1(n12784), .IN2(n12786), .QN(\fadd_0_0_0_0_9/newx [11])
         );
  NAND2X1 U6680 ( .IN1(n12737), .IN2(n12736), .QN(\fadd_0_0_0_0_4/newx [11])
         );
  NAND2X1 U6681 ( .IN1(n12757), .IN2(n12756), .QN(\fadd_0_0_0_0_6/newx [11])
         );
  NAND2X1 U6682 ( .IN1(n12764), .IN2(n12766), .QN(\fadd_0_0_0_0_7/newx [11])
         );
  NAND2X1 U6683 ( .IN1(n12744), .IN2(n12746), .QN(\fadd_0_0_0_0_5/newx [11])
         );
  NAND2X1 U6684 ( .IN1(n12717), .IN2(n12716), .QN(\fadd_0_0_0_0_2/newx [11])
         );
  NAND2X1 U6685 ( .IN1(n12724), .IN2(n12726), .QN(\fadd_0_0_0_0_3/newx [11])
         );
  NAND2X1 U6686 ( .IN1(n12704), .IN2(n12706), .QN(\fadd_0_0_0_0_1/newx [11])
         );
  XOR2X1 U6687 ( .IN1(n14171), .IN2(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/B[6] ), .Q(\fadd_0_0_0_0_10/U21/DATA2_3 ) );
  XOR2X1 U6688 ( .IN1(n14173), .IN2(
        \fmul_0_0_0_0_10/sub_1_root_add_321/carry[5] ), .Q(
        \fmul_0_0_0_0_10/sub_1_root_add_321/DIFF[5] ) );
  XOR2X1 U6689 ( .IN1(n14175), .IN2(n14122), .Q(
        \fmul_0_0_0_0_10/sub_1_root_add_321/DIFF[4] ) );
  XOR2X1 U6690 ( .IN1(n13467), .IN2(n14962), .Q(\fadd_0_0_0_0_10/U24/DATA2_1 )
         );
  XOR2X1 U6691 ( .IN1(n13884), .IN2(\fadd_0_0_0_0_10/sub_784/carry[4] ), .Q(
        \fadd_0_0_0_0_10/sub_784/DIFF[4] ) );
  XOR2X1 U6692 ( .IN1(n13749), .IN2(\fadd_0_0_0_0_10/sub_784/carry[3] ), .Q(
        \fadd_0_0_0_0_10/sub_784/DIFF[3] ) );
  XOR2X1 U6693 ( .IN1(n13714), .IN2(\fadd_0_0_0_0_10/norm/U5/Z_5 ), .Q(
        \fadd_0_0_0_0_10/sub_784/DIFF[0] ) );
  XOR2X1 U6694 ( .IN1(n14179), .IN2(n14180), .Q(\fadd_0_0_0_0_10/U5/DATA1_0 )
         );
  XOR2X1 U6695 ( .IN1(n14180), .IN2(n14179), .Q(\fadd_0_0_0_0_10/U5/DATA2_0 )
         );
  XOR2X1 U6696 ( .IN1(n14181), .IN2(\fadd_0_0_0_0_10/U27/DATA1_0 ), .Q(
        \fadd_0_0_0_0_10/U24/DATA1_5 ) );
  XOR2X1 U6697 ( .IN1(n14158), .IN2(
        \fmul_0_0_0_0_10/roundingadder/add_1_root_add_57/A[9] ), .Q(
        \fmul_0_0_0_0_10/roundingadder/add_1_root_add_57/SUM[9] ) );
  XOR2X1 U6698 ( .IN1(n14157), .IN2(
        \fmul_0_0_0_0_10/roundingadder/add_1_root_add_57/A[8] ), .Q(n13444) );
  XOR2X1 U6699 ( .IN1(n14160), .IN2(
        \fmul_0_0_0_0_10/roundingadder/add_1_root_add_57/A[7] ), .Q(n13445) );
  XOR2X1 U6700 ( .IN1(n14156), .IN2(
        \fmul_0_0_0_0_10/roundingadder/add_1_root_add_57/A[6] ), .Q(n13446) );
  XOR2X1 U6701 ( .IN1(n14155), .IN2(
        \fmul_0_0_0_0_10/roundingadder/add_1_root_add_57/A[5] ), .Q(n13447) );
  XOR2X1 U6702 ( .IN1(n14154), .IN2(
        \fmul_0_0_0_0_10/roundingadder/add_1_root_add_57/A[4] ), .Q(n13448) );
  XOR2X1 U6703 ( .IN1(n14153), .IN2(
        \fmul_0_0_0_0_10/roundingadder/add_1_root_add_57/A[3] ), .Q(n13449) );
  XOR2X1 U6704 ( .IN1(n14152), .IN2(
        \fmul_0_0_0_0_10/roundingadder/add_1_root_add_57/A[2] ), .Q(n13450) );
  XOR2X1 U6705 ( .IN1(n14151), .IN2(
        \fmul_0_0_0_0_10/roundingadder/add_1_root_add_57/A[1] ), .Q(n13451) );
  XOR2X1 U6706 ( .IN1(\fmul_0_0_0_0_10/roundingadder/add_1_root_add_57/CI ), 
        .IN2(\fmul_0_0_0_0_10/roundingadder/add_1_root_add_57/A[0] ), .Q(
        n13452) );
  XOR2X1 U6707 ( .IN1(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/B[7] ), .IN2(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/carry[7] ), .Q(\fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/SUM[7] ) );
  XOR2X1 U6708 ( .IN1(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/B[1] ), .IN2(n14139), .Q(\fadd_0_0_0_0_10/U22/DATA1_0 ) );
  XOR2X1 U6709 ( .IN1(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/B[0] ), .IN2(\fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_fracaddfar/add_1_root_add_54/CI ), 
        .Q(\fadd_0_0_0_0_10/U20/DATA1_0 ) );
  XOR2X1 U6710 ( .IN1(n13412), .IN2(\fadd_0_0_0_0_10/add_859/carry[6] ), .Q(
        \fadd_0_0_0_0_10/U4/DATA2_10 ) );
  XOR2X1 U6711 ( .IN1(n14121), .IN2(\fmul_0_0_0_0_10/sub_1_root_add_321/A[3] ), 
        .Q(\fmul_0_0_0_0_10/sub_1_root_add_321/DIFF[3] ) );
  XOR2X1 U6712 ( .IN1(n14120), .IN2(\fmul_0_0_0_0_10/sub_1_root_add_321/A[2] ), 
        .Q(\fmul_0_0_0_0_10/sub_1_root_add_321/DIFF[2] ) );
  XOR2X1 U6713 ( .IN1(\fmul_0_0_0_0_10/sub_1_root_add_321/A[0] ), .IN2(
        \fmul_0_0_0_0_10/sub_1_root_add_321/A[1] ), .Q(
        \fmul_0_0_0_0_10/sub_1_root_add_321/DIFF[1] ) );
  XOR2X1 U6714 ( .IN1(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_dualsubclose/sub_1_root_add_303/carry[5] ), .IN2(n14979), .Q(\fadd_0_0_0_0_10/U24/DATA2_5 ) );
  INVX0 U6715 ( .INP(n12829), .ZN(n14916) );
  INVX0 U6716 ( .INP(n12829), .ZN(n14201) );
  INVX0 U6717 ( .INP(n12829), .ZN(n14206) );
  INVX0 U6718 ( .INP(n12829), .ZN(n14202) );
  INVX0 U6719 ( .INP(n12829), .ZN(n14204) );
  INVX0 U6720 ( .INP(n12829), .ZN(n14205) );
  INVX0 U6721 ( .INP(n12829), .ZN(n14203) );
  INVX0 U6722 ( .INP(n12827), .ZN(n14184) );
  INVX0 U6723 ( .INP(n12827), .ZN(n14917) );
  INVX0 U6724 ( .INP(n11927), .ZN(n14914) );
  INVX0 U6725 ( .INP(n11927), .ZN(n14257) );
  INVX0 U6726 ( .INP(n11927), .ZN(n14256) );
  INVX0 U6727 ( .INP(n11927), .ZN(n14190) );
  INVX0 U6728 ( .INP(n11927), .ZN(n14193) );
  INVX0 U6729 ( .INP(n11927), .ZN(n14189) );
  INVX0 U6730 ( .INP(n11927), .ZN(n14191) );
  INVX0 U6731 ( .INP(n11927), .ZN(n14192) );
  AND2X1 U6732 ( .IN1(n8764), .IN2(n9130), .Q(n9166) );
  INVX0 U6733 ( .INP(n14435), .ZN(n14434) );
  INVX0 U6734 ( .INP(n14435), .ZN(n14209) );
  INVX0 U6735 ( .INP(n14435), .ZN(n14213) );
  INVX0 U6736 ( .INP(n14435), .ZN(n14214) );
  INVX0 U6737 ( .INP(n14435), .ZN(n14212) );
  INVX0 U6738 ( .INP(n14435), .ZN(n14207) );
  INVX0 U6739 ( .INP(n14435), .ZN(n14208) );
  INVX0 U6740 ( .INP(n14435), .ZN(n14210) );
  INVX0 U6741 ( .INP(n14435), .ZN(n14211) );
  INVX0 U6742 ( .INP(n11271), .ZN(n14188) );
  INVX0 U6743 ( .INP(n11271), .ZN(n14304) );
  INVX0 U6744 ( .INP(n10698), .ZN(n14311) );
  INVX0 U6745 ( .INP(n11105), .ZN(n14306) );
  INVX0 U6746 ( .INP(n10781), .ZN(n14310) );
  INVX0 U6747 ( .INP(n10617), .ZN(n14312) );
  INVX0 U6748 ( .INP(n10862), .ZN(n14309) );
  INVX0 U6749 ( .INP(n11322), .ZN(n14303) );
  INVX0 U6750 ( .INP(n11024), .ZN(n14307) );
  INVX0 U6751 ( .INP(n10943), .ZN(n14308) );
  INVX0 U6752 ( .INP(n11186), .ZN(n14305) );
  INVX0 U6753 ( .INP(n11403), .ZN(n14302) );
  NOR2X0 U6754 ( .IN1(n14437), .IN2(n12827), .QN(\U4/Z_44 ) );
  NOR2X0 U6755 ( .IN1(n14185), .IN2(n9057), .QN(n9129) );
  NBUFFX2 U6756 ( .INP(n9451), .Z(n14344) );
  INVX0 U6757 ( .INP(n14137), .ZN(n14436) );
  INVX0 U6758 ( .INP(n12828), .ZN(n14263) );
  NAND2X0 U6759 ( .IN1(n11241), .IN2(n11242), .QN(n11239) );
  INVX0 U6760 ( .INP(n14279), .ZN(n14277) );
  INVX0 U6761 ( .INP(n14279), .ZN(n14278) );
  INVX0 U6762 ( .INP(n14218), .ZN(n14220) );
  INVX0 U6763 ( .INP(n14218), .ZN(n14219) );
  INVX0 U6764 ( .INP(n12364), .ZN(n14282) );
  INVX0 U6765 ( .INP(n14281), .ZN(n14280) );
  INVX0 U6766 ( .INP(n14281), .ZN(n14279) );
  INVX0 U6767 ( .INP(n14277), .ZN(n14218) );
  INVX0 U6768 ( .INP(n14274), .ZN(n14272) );
  INVX0 U6769 ( .INP(n14274), .ZN(n14273) );
  INVX0 U6770 ( .INP(n14275), .ZN(n14269) );
  INVX0 U6771 ( .INP(n14275), .ZN(n14270) );
  INVX0 U6772 ( .INP(n14275), .ZN(n14271) );
  INVX0 U6773 ( .INP(n14276), .ZN(n14266) );
  INVX0 U6774 ( .INP(n14276), .ZN(n14267) );
  INVX0 U6775 ( .INP(n14276), .ZN(n14268) );
  INVX0 U6776 ( .INP(n14219), .ZN(n14265) );
  INVX0 U6777 ( .INP(n14219), .ZN(n14264) );
  INVX0 U6778 ( .INP(n14298), .ZN(n14296) );
  INVX0 U6779 ( .INP(n14298), .ZN(n14297) );
  INVX0 U6780 ( .INP(n14221), .ZN(n14223) );
  INVX0 U6781 ( .INP(n14221), .ZN(n14222) );
  INVX0 U6782 ( .INP(n12356), .ZN(n14301) );
  INVX0 U6783 ( .INP(n14300), .ZN(n14299) );
  INVX0 U6784 ( .INP(n14300), .ZN(n14298) );
  INVX0 U6785 ( .INP(n14296), .ZN(n14221) );
  INVX0 U6786 ( .INP(n14293), .ZN(n14291) );
  INVX0 U6787 ( .INP(n14293), .ZN(n14292) );
  INVX0 U6788 ( .INP(n14294), .ZN(n14288) );
  INVX0 U6789 ( .INP(n14294), .ZN(n14289) );
  INVX0 U6790 ( .INP(n14294), .ZN(n14290) );
  INVX0 U6791 ( .INP(n14295), .ZN(n14285) );
  INVX0 U6792 ( .INP(n14295), .ZN(n14286) );
  INVX0 U6793 ( .INP(n14295), .ZN(n14287) );
  INVX0 U6794 ( .INP(n14222), .ZN(n14284) );
  INVX0 U6795 ( .INP(n14222), .ZN(n14283) );
  INVX0 U6796 ( .INP(\fadd_0_0_0_0_10/U27/Z_2 ), .ZN(n14976) );
  NOR2X0 U6797 ( .IN1(\fadd_0_0_0_0_10/U27/Z_1 ), .IN2(
        \fadd_0_0_0_0_10/U27/Z_2 ), .QN(n11241) );
  NAND2X0 U6798 ( .IN1(\fadd_0_0_0_0_10/U27/Z_2 ), .IN2(n14974), .QN(n11234)
         );
  NOR2X0 U6799 ( .IN1(n14965), .IN2(\fadd_0_0_0_0_10/U27/Z_2 ), .QN(n11258) );
  OA22X1 U6800 ( .IN1(n11284), .IN2(n12808), .IN3(n13500), .IN4(n11285), .Q(
        n11271) );
  INVX0 U6801 ( .INP(n8766), .ZN(n14435) );
  NOR2X0 U6802 ( .IN1(n14183), .IN2(n14187), .QN(n8764) );
  NAND2X0 U6803 ( .IN1(n14113), .IN2(n14672), .QN(n11315) );
  NAND2X0 U6804 ( .IN1(n14117), .IN2(n14725), .QN(n11098) );
  NAND2X0 U6805 ( .IN1(n14111), .IN2(n14778), .QN(n10936) );
  NAND2X0 U6806 ( .IN1(n14116), .IN2(n14820), .QN(n10774) );
  NAND2X0 U6807 ( .IN1(n14110), .IN2(n14746), .QN(n11017) );
  NAND2X0 U6808 ( .IN1(n14114), .IN2(n14873), .QN(n10610) );
  NAND2X0 U6809 ( .IN1(n14112), .IN2(n14693), .QN(n11179) );
  NAND2X0 U6810 ( .IN1(n14115), .IN2(n14799), .QN(n10855) );
  NAND2X0 U6811 ( .IN1(n14109), .IN2(n14651), .QN(n11396) );
  NAND2X0 U6812 ( .IN1(n14118), .IN2(n14841), .QN(n10691) );
  INVX0 U6813 ( .INP(
        \fadd_0_0_0_0_10/fpadd_5_4_f300_uid2_dualsubclose/sub_1_root_add_300/carry[6] ), .ZN(n14963) );
  NOR2X0 U6814 ( .IN1(n8990), .IN2(n9097), .QN(n9410) );
  NOR2X0 U6815 ( .IN1(n9130), .IN2(n14185), .QN(n9057) );
  INVX0 U6816 ( .INP(n9057), .ZN(n14419) );
  XNOR2X1 U6817 ( .IN1(\fadd_0_0_0_0_8/newx_d1 [8]), .IN2(
        \fadd_0_0_0_0_8/sub_784/carry [4]), .Q(
        \fadd_0_0_0_0_8/exponentresultclose [4]) );
  OR2X1 U6818 ( .IN1(\fadd_0_0_0_0_8/sub_784/carry [3]), .IN2(
        \fadd_0_0_0_0_8/newx_d1 [7]), .Q(\fadd_0_0_0_0_8/sub_784/carry [4]) );
  XNOR2X1 U6819 ( .IN1(\fadd_0_0_0_0_8/newx_d1 [7]), .IN2(
        \fadd_0_0_0_0_8/sub_784/carry [3]), .Q(
        \fadd_0_0_0_0_8/exponentresultclose [3]) );
  OR2X1 U6820 ( .IN1(n14629), .IN2(\fadd_0_0_0_0_8/newx_d1 [4]), .Q(
        \fadd_0_0_0_0_8/sub_784/carry [1]) );
  XNOR2X1 U6821 ( .IN1(\fadd_0_0_0_0_8/newx_d1 [4]), .IN2(n14629), .Q(
        \fadd_0_0_0_0_8/exponentresultclose [0]) );
  XOR2X1 U6822 ( .IN1(
        \add_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [10]), .IN2(\fadd_0_0_0_0_8/resultbeforeround [10]), .Q(
        \fadd_0_0_0_0_8/resultrounded [10]) );
  XOR2X1 U6823 ( .IN1(\fadd_0_0_0_0_8/add_859/B[1] ), .IN2(
        \fadd_0_0_0_0_8/add_859/carry [6]), .Q(
        \fadd_0_0_0_0_8/exponentresultfar1 [6]) );
  AND2X1 U6824 ( .IN1(
        \add_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [9]), .IN2(\fadd_0_0_0_0_8/resultbeforeround [9]), .Q(
        \add_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [10]) );
  AND2X1 U6825 ( .IN1(
        \add_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [8]), .IN2(\fadd_0_0_0_0_8/resultbeforeround [8]), .Q(
        \add_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [9]) );
  XOR2X1 U6826 ( .IN1(
        \add_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [8]), .IN2(\fadd_0_0_0_0_8/resultbeforeround [8]), .Q(
        \fadd_0_0_0_0_8/resultrounded [8]) );
  AND2X1 U6827 ( .IN1(
        \add_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [7]), .IN2(\fadd_0_0_0_0_8/resultbeforeround [7]), .Q(
        \add_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [8]) );
  XOR2X1 U6828 ( .IN1(
        \add_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [7]), .IN2(\fadd_0_0_0_0_8/resultbeforeround [7]), .Q(
        \fadd_0_0_0_0_8/resultrounded [7]) );
  AND2X1 U6829 ( .IN1(
        \add_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [6]), .IN2(\fadd_0_0_0_0_8/resultbeforeround [6]), .Q(
        \add_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [7]) );
  XOR2X1 U6830 ( .IN1(
        \add_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [6]), .IN2(\fadd_0_0_0_0_8/resultbeforeround [6]), .Q(
        \fadd_0_0_0_0_8/resultrounded [6]) );
  AND2X1 U6831 ( .IN1(
        \add_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [5]), .IN2(\fadd_0_0_0_0_8/resultbeforeround [5]), .Q(
        \add_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [6]) );
  XOR2X1 U6832 ( .IN1(
        \add_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [5]), .IN2(\fadd_0_0_0_0_8/resultbeforeround [5]), .Q(
        \fadd_0_0_0_0_8/resultrounded [5]) );
  AND2X1 U6833 ( .IN1(
        \add_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [4]), .IN2(\fadd_0_0_0_0_8/resultbeforeround [4]), .Q(
        \add_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [5]) );
  XOR2X1 U6834 ( .IN1(
        \add_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [4]), .IN2(\fadd_0_0_0_0_8/resultbeforeround [4]), .Q(
        \fadd_0_0_0_0_8/resultrounded [4]) );
  AND2X1 U6835 ( .IN1(
        \add_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [3]), .IN2(\fadd_0_0_0_0_8/resultbeforeround [3]), .Q(
        \add_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [4]) );
  XOR2X1 U6836 ( .IN1(
        \add_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [3]), .IN2(\fadd_0_0_0_0_8/resultbeforeround [3]), .Q(
        \fadd_0_0_0_0_8/resultrounded [3]) );
  AND2X1 U6837 ( .IN1(
        \add_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [2]), .IN2(\fadd_0_0_0_0_8/resultbeforeround [2]), .Q(
        \add_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [3]) );
  XOR2X1 U6838 ( .IN1(
        \add_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [2]), .IN2(\fadd_0_0_0_0_8/resultbeforeround [2]), .Q(
        \fadd_0_0_0_0_8/resultrounded [2]) );
  AND2X1 U6839 ( .IN1(
        \add_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [1]), .IN2(\fadd_0_0_0_0_8/resultbeforeround [1]), .Q(
        \add_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [2]) );
  XOR2X1 U6840 ( .IN1(
        \add_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [1]), .IN2(\fadd_0_0_0_0_8/resultbeforeround [1]), .Q(
        \fadd_0_0_0_0_8/resultrounded [1]) );
  AND2X1 U6841 ( .IN1(\fadd_0_0_0_0_8/round ), .IN2(
        \fadd_0_0_0_0_8/resultbeforeround [0]), .Q(
        \add_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [1]) );
  XOR2X1 U6842 ( .IN1(\fadd_0_0_0_0_8/round ), .IN2(
        \fadd_0_0_0_0_8/resultbeforeround [0]), .Q(
        \fadd_0_0_0_0_8/resultrounded [0]) );
  AND2X1 U6843 ( .IN1(\fadd_0_0_0_0_8/add_859/B[1] ), .IN2(
        \fadd_0_0_0_0_8/add_859/carry [5]), .Q(
        \fadd_0_0_0_0_8/add_859/carry [6]) );
  XOR2X1 U6844 ( .IN1(\fadd_0_0_0_0_8/add_859/B[1] ), .IN2(
        \fadd_0_0_0_0_8/add_859/carry [5]), .Q(
        \fadd_0_0_0_0_8/exponentresultfar1 [5]) );
  AND2X1 U6845 ( .IN1(\fadd_0_0_0_0_8/expoperationsel[0] ), .IN2(
        \fadd_0_0_0_0_8/exponentresultfar0_d2 [0]), .Q(
        \fadd_0_0_0_0_8/add_859/carry [1]) );
  XOR2X1 U6846 ( .IN1(\fadd_0_0_0_0_8/expoperationsel[0] ), .IN2(
        \fadd_0_0_0_0_8/exponentresultfar0_d2 [0]), .Q(
        \fadd_0_0_0_0_8/exponentresultfar1 [0]) );
  XOR2X1 U6847 ( .IN1(
        \add_1_root_fmul_0_0_0_0_8/roundingadder/add_57/carry [10]), .IN2(
        \fmul_0_0_0_0_8/roundingadder/x_1_d1 [10]), .Q(
        \fmul_0_0_0_0_8/expsigpostround[10] ) );
  AND2X1 U6848 ( .IN1(
        \add_1_root_fmul_0_0_0_0_8/roundingadder/add_57/carry [9]), .IN2(
        \fmul_0_0_0_0_8/roundingadder/x_1_d1 [9]), .Q(
        \add_1_root_fmul_0_0_0_0_8/roundingadder/add_57/carry [10]) );
  AND2X1 U6849 ( .IN1(\fmul_0_0_0_0_8/roundingadder/x_1_d1 [8]), .IN2(
        \add_1_root_fmul_0_0_0_0_8/roundingadder/add_57/carry [8]), .Q(
        \add_1_root_fmul_0_0_0_0_8/roundingadder/add_57/carry [9]) );
  XOR2X1 U6850 ( .IN1(
        \add_1_root_fmul_0_0_0_0_8/roundingadder/add_57/carry [8]), .IN2(
        \fmul_0_0_0_0_8/roundingadder/x_1_d1 [8]), .Q(\U120/DATA2_8 ) );
  AND2X1 U6851 ( .IN1(\fmul_0_0_0_0_8/roundingadder/x_1_d1 [7]), .IN2(
        \add_1_root_fmul_0_0_0_0_8/roundingadder/add_57/carry [7]), .Q(
        \add_1_root_fmul_0_0_0_0_8/roundingadder/add_57/carry [8]) );
  XOR2X1 U6852 ( .IN1(
        \add_1_root_fmul_0_0_0_0_8/roundingadder/add_57/carry [7]), .IN2(
        \fmul_0_0_0_0_8/roundingadder/x_1_d1 [7]), .Q(\U120/DATA2_7 ) );
  AND2X1 U6853 ( .IN1(\fmul_0_0_0_0_8/roundingadder/x_1_d1 [6]), .IN2(
        \add_1_root_fmul_0_0_0_0_8/roundingadder/add_57/carry [6]), .Q(
        \add_1_root_fmul_0_0_0_0_8/roundingadder/add_57/carry [7]) );
  XOR2X1 U6854 ( .IN1(
        \add_1_root_fmul_0_0_0_0_8/roundingadder/add_57/carry [6]), .IN2(
        \fmul_0_0_0_0_8/roundingadder/x_1_d1 [6]), .Q(\U120/DATA2_6 ) );
  AND2X1 U6855 ( .IN1(\fmul_0_0_0_0_8/roundingadder/x_1_d1 [5]), .IN2(
        \add_1_root_fmul_0_0_0_0_8/roundingadder/add_57/carry [5]), .Q(
        \add_1_root_fmul_0_0_0_0_8/roundingadder/add_57/carry [6]) );
  XOR2X1 U6856 ( .IN1(
        \add_1_root_fmul_0_0_0_0_8/roundingadder/add_57/carry [5]), .IN2(
        \fmul_0_0_0_0_8/roundingadder/x_1_d1 [5]), .Q(\U120/DATA2_5 ) );
  AND2X1 U6857 ( .IN1(\fmul_0_0_0_0_8/roundingadder/x_1_d1 [4]), .IN2(
        \add_1_root_fmul_0_0_0_0_8/roundingadder/add_57/carry [4]), .Q(
        \add_1_root_fmul_0_0_0_0_8/roundingadder/add_57/carry [5]) );
  XOR2X1 U6858 ( .IN1(
        \add_1_root_fmul_0_0_0_0_8/roundingadder/add_57/carry [4]), .IN2(
        \fmul_0_0_0_0_8/roundingadder/x_1_d1 [4]), .Q(\U120/DATA2_4 ) );
  AND2X1 U6859 ( .IN1(\fmul_0_0_0_0_8/roundingadder/x_1_d1 [3]), .IN2(
        \add_1_root_fmul_0_0_0_0_8/roundingadder/add_57/carry [3]), .Q(
        \add_1_root_fmul_0_0_0_0_8/roundingadder/add_57/carry [4]) );
  XOR2X1 U6860 ( .IN1(
        \add_1_root_fmul_0_0_0_0_8/roundingadder/add_57/carry [3]), .IN2(
        \fmul_0_0_0_0_8/roundingadder/x_1_d1 [3]), .Q(\U120/DATA2_3 ) );
  AND2X1 U6861 ( .IN1(\fmul_0_0_0_0_8/roundingadder/x_1_d1 [2]), .IN2(
        \add_1_root_fmul_0_0_0_0_8/roundingadder/add_57/carry [2]), .Q(
        \add_1_root_fmul_0_0_0_0_8/roundingadder/add_57/carry [3]) );
  XOR2X1 U6862 ( .IN1(
        \add_1_root_fmul_0_0_0_0_8/roundingadder/add_57/carry [2]), .IN2(
        \fmul_0_0_0_0_8/roundingadder/x_1_d1 [2]), .Q(\U120/DATA2_2 ) );
  AND2X1 U6863 ( .IN1(\fmul_0_0_0_0_8/roundingadder/x_1_d1 [1]), .IN2(
        \add_1_root_fmul_0_0_0_0_8/roundingadder/add_57/carry [1]), .Q(
        \add_1_root_fmul_0_0_0_0_8/roundingadder/add_57/carry [2]) );
  XOR2X1 U6864 ( .IN1(
        \add_1_root_fmul_0_0_0_0_8/roundingadder/add_57/carry [1]), .IN2(
        \fmul_0_0_0_0_8/roundingadder/x_1_d1 [1]), .Q(\U120/DATA2_1 ) );
  AND2X1 U6865 ( .IN1(\fmul_0_0_0_0_8/roundingadder/x_1_d1 [0]), .IN2(
        \fmul_0_0_0_0_8/roundingadder/n151_o[0] ), .Q(
        \add_1_root_fmul_0_0_0_0_8/roundingadder/add_57/carry [1]) );
  XOR2X1 U6866 ( .IN1(\fmul_0_0_0_0_8/roundingadder/n151_o[0] ), .IN2(
        \fmul_0_0_0_0_8/roundingadder/x_1_d1 [0]), .Q(\U120/DATA2_0 ) );
  XNOR2X1 U6867 ( .IN1(\fadd_0_0_0_0_9/newx_d1 [8]), .IN2(
        \fadd_0_0_0_0_9/sub_784/carry [4]), .Q(
        \fadd_0_0_0_0_9/exponentresultclose [4]) );
  OR2X1 U6868 ( .IN1(\fadd_0_0_0_0_9/sub_784/carry [3]), .IN2(
        \fadd_0_0_0_0_9/newx_d1 [7]), .Q(\fadd_0_0_0_0_9/sub_784/carry [4]) );
  XNOR2X1 U6869 ( .IN1(\fadd_0_0_0_0_9/newx_d1 [7]), .IN2(
        \fadd_0_0_0_0_9/sub_784/carry [3]), .Q(
        \fadd_0_0_0_0_9/exponentresultclose [3]) );
  OR2X1 U6870 ( .IN1(n14640), .IN2(\fadd_0_0_0_0_9/newx_d1 [4]), .Q(
        \fadd_0_0_0_0_9/sub_784/carry [1]) );
  XNOR2X1 U6871 ( .IN1(\fadd_0_0_0_0_9/newx_d1 [4]), .IN2(n14640), .Q(
        \fadd_0_0_0_0_9/exponentresultclose [0]) );
  XOR2X1 U6872 ( .IN1(
        \add_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [10]), .IN2(\fadd_0_0_0_0_9/resultbeforeround [10]), .Q(
        \fadd_0_0_0_0_9/resultrounded [10]) );
  XOR2X1 U6873 ( .IN1(\fadd_0_0_0_0_9/add_859/B[1] ), .IN2(
        \fadd_0_0_0_0_9/add_859/carry [6]), .Q(
        \fadd_0_0_0_0_9/exponentresultfar1 [6]) );
  AND2X1 U6874 ( .IN1(
        \add_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [9]), .IN2(\fadd_0_0_0_0_9/resultbeforeround [9]), .Q(
        \add_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [10]) );
  XOR2X1 U6875 ( .IN1(
        \add_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [9]), .IN2(\fadd_0_0_0_0_9/resultbeforeround [9]), .Q(
        \fadd_0_0_0_0_9/resultrounded [9]) );
  AND2X1 U6876 ( .IN1(
        \add_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [8]), .IN2(\fadd_0_0_0_0_9/resultbeforeround [8]), .Q(
        \add_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [9]) );
  XOR2X1 U6877 ( .IN1(
        \add_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [8]), .IN2(\fadd_0_0_0_0_9/resultbeforeround [8]), .Q(
        \fadd_0_0_0_0_9/resultrounded [8]) );
  AND2X1 U6878 ( .IN1(
        \add_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [7]), .IN2(\fadd_0_0_0_0_9/resultbeforeround [7]), .Q(
        \add_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [8]) );
  XOR2X1 U6879 ( .IN1(
        \add_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [7]), .IN2(\fadd_0_0_0_0_9/resultbeforeround [7]), .Q(
        \fadd_0_0_0_0_9/resultrounded [7]) );
  AND2X1 U6880 ( .IN1(
        \add_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [6]), .IN2(\fadd_0_0_0_0_9/resultbeforeround [6]), .Q(
        \add_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [7]) );
  XOR2X1 U6881 ( .IN1(
        \add_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [6]), .IN2(\fadd_0_0_0_0_9/resultbeforeround [6]), .Q(
        \fadd_0_0_0_0_9/resultrounded [6]) );
  AND2X1 U6882 ( .IN1(
        \add_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [5]), .IN2(\fadd_0_0_0_0_9/resultbeforeround [5]), .Q(
        \add_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [6]) );
  XOR2X1 U6883 ( .IN1(
        \add_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [5]), .IN2(\fadd_0_0_0_0_9/resultbeforeround [5]), .Q(
        \fadd_0_0_0_0_9/resultrounded [5]) );
  AND2X1 U6884 ( .IN1(
        \add_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [4]), .IN2(\fadd_0_0_0_0_9/resultbeforeround [4]), .Q(
        \add_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [5]) );
  XOR2X1 U6885 ( .IN1(
        \add_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [4]), .IN2(\fadd_0_0_0_0_9/resultbeforeround [4]), .Q(
        \fadd_0_0_0_0_9/resultrounded [4]) );
  AND2X1 U6886 ( .IN1(
        \add_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [3]), .IN2(\fadd_0_0_0_0_9/resultbeforeround [3]), .Q(
        \add_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [4]) );
  XOR2X1 U6887 ( .IN1(
        \add_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [3]), .IN2(\fadd_0_0_0_0_9/resultbeforeround [3]), .Q(
        \fadd_0_0_0_0_9/resultrounded [3]) );
  AND2X1 U6888 ( .IN1(
        \add_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [2]), .IN2(\fadd_0_0_0_0_9/resultbeforeround [2]), .Q(
        \add_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [3]) );
  XOR2X1 U6889 ( .IN1(
        \add_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [2]), .IN2(\fadd_0_0_0_0_9/resultbeforeround [2]), .Q(
        \fadd_0_0_0_0_9/resultrounded [2]) );
  AND2X1 U6890 ( .IN1(
        \add_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [1]), .IN2(\fadd_0_0_0_0_9/resultbeforeround [1]), .Q(
        \add_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [2]) );
  XOR2X1 U6891 ( .IN1(
        \add_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [1]), .IN2(\fadd_0_0_0_0_9/resultbeforeround [1]), .Q(
        \fadd_0_0_0_0_9/resultrounded [1]) );
  AND2X1 U6892 ( .IN1(\fadd_0_0_0_0_9/round ), .IN2(
        \fadd_0_0_0_0_9/resultbeforeround [0]), .Q(
        \add_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [1]) );
  XOR2X1 U6893 ( .IN1(\fadd_0_0_0_0_9/round ), .IN2(
        \fadd_0_0_0_0_9/resultbeforeround [0]), .Q(
        \fadd_0_0_0_0_9/resultrounded [0]) );
  AND2X1 U6894 ( .IN1(\fadd_0_0_0_0_9/add_859/B[1] ), .IN2(
        \fadd_0_0_0_0_9/add_859/carry [5]), .Q(
        \fadd_0_0_0_0_9/add_859/carry [6]) );
  XOR2X1 U6895 ( .IN1(\fadd_0_0_0_0_9/add_859/B[1] ), .IN2(
        \fadd_0_0_0_0_9/add_859/carry [5]), .Q(
        \fadd_0_0_0_0_9/exponentresultfar1 [5]) );
  AND2X1 U6896 ( .IN1(\fadd_0_0_0_0_9/expoperationsel[0] ), .IN2(
        \fadd_0_0_0_0_9/exponentresultfar0_d2 [0]), .Q(
        \fadd_0_0_0_0_9/add_859/carry [1]) );
  XOR2X1 U6897 ( .IN1(\fadd_0_0_0_0_9/expoperationsel[0] ), .IN2(
        \fadd_0_0_0_0_9/exponentresultfar0_d2 [0]), .Q(
        \fadd_0_0_0_0_9/exponentresultfar1 [0]) );
  XOR2X1 U6898 ( .IN1(
        \add_1_root_fmul_0_0_0_0_9/roundingadder/add_57/carry [10]), .IN2(
        \fmul_0_0_0_0_9/roundingadder/x_1_d1 [10]), .Q(
        \fmul_0_0_0_0_9/expsigpostround [10]) );
  AND2X1 U6899 ( .IN1(
        \add_1_root_fmul_0_0_0_0_9/roundingadder/add_57/carry [9]), .IN2(
        \fmul_0_0_0_0_9/roundingadder/x_1_d1 [9]), .Q(
        \add_1_root_fmul_0_0_0_0_9/roundingadder/add_57/carry [10]) );
  XOR2X1 U6900 ( .IN1(
        \add_1_root_fmul_0_0_0_0_9/roundingadder/add_57/carry [9]), .IN2(
        \fmul_0_0_0_0_9/roundingadder/x_1_d1 [9]), .Q(
        \fmul_0_0_0_0_9/expsigpostround [9]) );
  AND2X1 U6901 ( .IN1(\fmul_0_0_0_0_9/roundingadder/x_1_d1 [8]), .IN2(
        \add_1_root_fmul_0_0_0_0_9/roundingadder/add_57/carry [8]), .Q(
        \add_1_root_fmul_0_0_0_0_9/roundingadder/add_57/carry [9]) );
  XOR2X1 U6902 ( .IN1(
        \add_1_root_fmul_0_0_0_0_9/roundingadder/add_57/carry [8]), .IN2(
        \fmul_0_0_0_0_9/roundingadder/x_1_d1 [8]), .Q(\U58/DATA2_8 ) );
  AND2X1 U6903 ( .IN1(\fmul_0_0_0_0_9/roundingadder/x_1_d1 [7]), .IN2(
        \add_1_root_fmul_0_0_0_0_9/roundingadder/add_57/carry [7]), .Q(
        \add_1_root_fmul_0_0_0_0_9/roundingadder/add_57/carry [8]) );
  XOR2X1 U6904 ( .IN1(
        \add_1_root_fmul_0_0_0_0_9/roundingadder/add_57/carry [7]), .IN2(
        \fmul_0_0_0_0_9/roundingadder/x_1_d1 [7]), .Q(\U58/DATA2_7 ) );
  AND2X1 U6905 ( .IN1(\fmul_0_0_0_0_9/roundingadder/x_1_d1 [6]), .IN2(
        \add_1_root_fmul_0_0_0_0_9/roundingadder/add_57/carry [6]), .Q(
        \add_1_root_fmul_0_0_0_0_9/roundingadder/add_57/carry [7]) );
  XOR2X1 U6906 ( .IN1(
        \add_1_root_fmul_0_0_0_0_9/roundingadder/add_57/carry [6]), .IN2(
        \fmul_0_0_0_0_9/roundingadder/x_1_d1 [6]), .Q(\U58/DATA2_6 ) );
  AND2X1 U6907 ( .IN1(\fmul_0_0_0_0_9/roundingadder/x_1_d1 [5]), .IN2(
        \add_1_root_fmul_0_0_0_0_9/roundingadder/add_57/carry [5]), .Q(
        \add_1_root_fmul_0_0_0_0_9/roundingadder/add_57/carry [6]) );
  XOR2X1 U6908 ( .IN1(
        \add_1_root_fmul_0_0_0_0_9/roundingadder/add_57/carry [5]), .IN2(
        \fmul_0_0_0_0_9/roundingadder/x_1_d1 [5]), .Q(\U58/DATA2_5 ) );
  AND2X1 U6909 ( .IN1(\fmul_0_0_0_0_9/roundingadder/x_1_d1 [4]), .IN2(
        \add_1_root_fmul_0_0_0_0_9/roundingadder/add_57/carry [4]), .Q(
        \add_1_root_fmul_0_0_0_0_9/roundingadder/add_57/carry [5]) );
  XOR2X1 U6910 ( .IN1(
        \add_1_root_fmul_0_0_0_0_9/roundingadder/add_57/carry [4]), .IN2(
        \fmul_0_0_0_0_9/roundingadder/x_1_d1 [4]), .Q(\U58/DATA2_4 ) );
  AND2X1 U6911 ( .IN1(
        \add_1_root_fmul_0_0_0_0_9/roundingadder/add_57/carry [3]), .IN2(
        \fmul_0_0_0_0_9/roundingadder/x_1_d1 [3]), .Q(
        \add_1_root_fmul_0_0_0_0_9/roundingadder/add_57/carry [4]) );
  XOR2X1 U6912 ( .IN1(
        \add_1_root_fmul_0_0_0_0_9/roundingadder/add_57/carry [3]), .IN2(
        \fmul_0_0_0_0_9/roundingadder/x_1_d1 [3]), .Q(n13453) );
  AND2X1 U6913 ( .IN1(
        \add_1_root_fmul_0_0_0_0_9/roundingadder/add_57/carry [2]), .IN2(
        \fmul_0_0_0_0_9/roundingadder/x_1_d1 [2]), .Q(
        \add_1_root_fmul_0_0_0_0_9/roundingadder/add_57/carry [3]) );
  XOR2X1 U6914 ( .IN1(
        \add_1_root_fmul_0_0_0_0_9/roundingadder/add_57/carry [2]), .IN2(
        \fmul_0_0_0_0_9/roundingadder/x_1_d1 [2]), .Q(n13454) );
  AND2X1 U6915 ( .IN1(
        \add_1_root_fmul_0_0_0_0_9/roundingadder/add_57/carry [1]), .IN2(
        \fmul_0_0_0_0_9/roundingadder/x_1_d1 [1]), .Q(
        \add_1_root_fmul_0_0_0_0_9/roundingadder/add_57/carry [2]) );
  XOR2X1 U6916 ( .IN1(
        \add_1_root_fmul_0_0_0_0_9/roundingadder/add_57/carry [1]), .IN2(
        \fmul_0_0_0_0_9/roundingadder/x_1_d1 [1]), .Q(n13455) );
  AND2X1 U6917 ( .IN1(\fmul_0_0_0_0_9/roundingadder/n151_o[0] ), .IN2(
        \fmul_0_0_0_0_9/roundingadder/x_1_d1 [0]), .Q(
        \add_1_root_fmul_0_0_0_0_9/roundingadder/add_57/carry [1]) );
  XOR2X1 U6918 ( .IN1(\fmul_0_0_0_0_9/roundingadder/n151_o[0] ), .IN2(
        \fmul_0_0_0_0_9/roundingadder/x_1_d1 [0]), .Q(n13456) );
  XNOR2X1 U6919 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/A[5] ), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/carry [5]), .Q(
        \fmul_0_0_0_0_9/exppostnorm [5]) );
  OR2X1 U6920 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/carry [4]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/A[4] ), .Q(
        \add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/carry [5]) );
  XNOR2X1 U6921 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/A[4] ), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/carry [4]), .Q(
        \fmul_0_0_0_0_9/exppostnorm [4]) );
  AND2X1 U6922 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/carry [3]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/A[3] ), .Q(
        \add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/carry [4]) );
  XOR2X1 U6923 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/carry [3]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/A[3] ), .Q(
        \fmul_0_0_0_0_9/exppostnorm [3]) );
  AND2X1 U6924 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/carry [2]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/A[2] ), .Q(
        \add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/carry [3]) );
  XOR2X1 U6925 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/carry [2]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/A[2] ), .Q(
        \fmul_0_0_0_0_9/exppostnorm [2]) );
  AND2X1 U6926 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/B[0] ), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/A[0] ), .Q(
        \add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/carry [1]) );
  XOR2X1 U6927 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/B[0] ), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/A[0] ), .Q(
        \fmul_0_0_0_0_9/exppostnorm [0]) );
  AND2X1 U6928 ( .IN1(n5310), .IN2(n5298), .Q(
        \add_2_root_sub_1_root_fmul_0_0_0_0_9/add_321/carry [1]) );
  XOR2X1 U6929 ( .IN1(n5298), .IN2(n5310), .Q(
        \add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/A[0] ) );
  XNOR2X1 U6930 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/A[5] ), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/carry [5]), .Q(
        \fmul_0_0_0_0_8/exppostnorm [5]) );
  OR2X1 U6931 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/carry [4]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/A[4] ), .Q(
        \add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/carry [5]) );
  XNOR2X1 U6932 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/A[4] ), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/carry [4]), .Q(
        \fmul_0_0_0_0_8/exppostnorm [4]) );
  AND2X1 U6933 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/carry [3]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/A[3] ), .Q(
        \add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/carry [4]) );
  XOR2X1 U6934 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/carry [3]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/A[3] ), .Q(
        \fmul_0_0_0_0_8/exppostnorm [3]) );
  AND2X1 U6935 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/carry [2]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/A[2] ), .Q(
        \add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/carry [3]) );
  XOR2X1 U6936 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/carry [2]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/A[2] ), .Q(
        \fmul_0_0_0_0_8/exppostnorm [2]) );
  AND2X1 U6937 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/B[0] ), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/A[0] ), .Q(
        \add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/carry [1]) );
  XOR2X1 U6938 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/B[0] ), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/A[0] ), .Q(
        \fmul_0_0_0_0_8/exppostnorm [0]) );
  AND2X1 U6939 ( .IN1(n5382), .IN2(n5370), .Q(
        \add_2_root_sub_1_root_fmul_0_0_0_0_8/add_321/carry [1]) );
  XOR2X1 U6940 ( .IN1(n5370), .IN2(n5382), .Q(
        \add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/A[0] ) );
  XNOR2X1 U6941 ( .IN1(\fadd_0_0_0_0_0/newx_d1 [8]), .IN2(
        \fadd_0_0_0_0_0/sub_784/carry [4]), .Q(
        \fadd_0_0_0_0_0/exponentresultclose [4]) );
  OR2X1 U6942 ( .IN1(\fadd_0_0_0_0_0/sub_784/carry [3]), .IN2(
        \fadd_0_0_0_0_0/newx_d1 [7]), .Q(\fadd_0_0_0_0_0/sub_784/carry [4]) );
  XNOR2X1 U6943 ( .IN1(\fadd_0_0_0_0_0/newx_d1 [7]), .IN2(
        \fadd_0_0_0_0_0/sub_784/carry [3]), .Q(
        \fadd_0_0_0_0_0/exponentresultclose [3]) );
  OR2X1 U6944 ( .IN1(n14541), .IN2(\fadd_0_0_0_0_0/newx_d1 [4]), .Q(
        \fadd_0_0_0_0_0/sub_784/carry [1]) );
  XNOR2X1 U6945 ( .IN1(\fadd_0_0_0_0_0/newx_d1 [4]), .IN2(n14541), .Q(
        \fadd_0_0_0_0_0/exponentresultclose [0]) );
  XOR2X1 U6946 ( .IN1(
        \add_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [10]), .IN2(\fadd_0_0_0_0_0/resultbeforeround [10]), .Q(
        \fadd_0_0_0_0_0/resultrounded [10]) );
  XOR2X1 U6947 ( .IN1(n14224), .IN2(\fadd_0_0_0_0_0/add_859/carry [6]), .Q(
        \fadd_0_0_0_0_0/exponentresultfar1 [6]) );
  AND2X1 U6948 ( .IN1(
        \add_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [9]), .IN2(\fadd_0_0_0_0_0/resultbeforeround [9]), .Q(
        \add_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [10]) );
  XOR2X1 U6949 ( .IN1(
        \add_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [9]), .IN2(\fadd_0_0_0_0_0/resultbeforeround [9]), .Q(
        \fadd_0_0_0_0_0/resultrounded [9]) );
  AND2X1 U6950 ( .IN1(
        \add_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [8]), .IN2(\fadd_0_0_0_0_0/resultbeforeround [8]), .Q(
        \add_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [9]) );
  XOR2X1 U6951 ( .IN1(
        \add_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [8]), .IN2(\fadd_0_0_0_0_0/resultbeforeround [8]), .Q(
        \fadd_0_0_0_0_0/resultrounded [8]) );
  AND2X1 U6952 ( .IN1(
        \add_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [7]), .IN2(\fadd_0_0_0_0_0/resultbeforeround [7]), .Q(
        \add_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [8]) );
  XOR2X1 U6953 ( .IN1(
        \add_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [7]), .IN2(\fadd_0_0_0_0_0/resultbeforeround [7]), .Q(
        \fadd_0_0_0_0_0/resultrounded [7]) );
  AND2X1 U6954 ( .IN1(
        \add_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [6]), .IN2(\fadd_0_0_0_0_0/resultbeforeround [6]), .Q(
        \add_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [7]) );
  XOR2X1 U6955 ( .IN1(
        \add_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [6]), .IN2(\fadd_0_0_0_0_0/resultbeforeround [6]), .Q(
        \fadd_0_0_0_0_0/resultrounded [6]) );
  AND2X1 U6956 ( .IN1(
        \add_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [5]), .IN2(\fadd_0_0_0_0_0/resultbeforeround [5]), .Q(
        \add_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [6]) );
  XOR2X1 U6957 ( .IN1(
        \add_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [5]), .IN2(\fadd_0_0_0_0_0/resultbeforeround [5]), .Q(
        \fadd_0_0_0_0_0/resultrounded [5]) );
  AND2X1 U6958 ( .IN1(
        \add_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [4]), .IN2(\fadd_0_0_0_0_0/resultbeforeround [4]), .Q(
        \add_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [5]) );
  XOR2X1 U6959 ( .IN1(
        \add_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [4]), .IN2(\fadd_0_0_0_0_0/resultbeforeround [4]), .Q(
        \fadd_0_0_0_0_0/resultrounded [4]) );
  AND2X1 U6960 ( .IN1(
        \add_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [3]), .IN2(\fadd_0_0_0_0_0/resultbeforeround [3]), .Q(
        \add_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [4]) );
  XOR2X1 U6961 ( .IN1(
        \add_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [3]), .IN2(\fadd_0_0_0_0_0/resultbeforeround [3]), .Q(
        \fadd_0_0_0_0_0/resultrounded [3]) );
  AND2X1 U6962 ( .IN1(
        \add_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [2]), .IN2(\fadd_0_0_0_0_0/resultbeforeround [2]), .Q(
        \add_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [3]) );
  XOR2X1 U6963 ( .IN1(
        \add_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [2]), .IN2(\fadd_0_0_0_0_0/resultbeforeround [2]), .Q(
        \fadd_0_0_0_0_0/resultrounded [2]) );
  AND2X1 U6964 ( .IN1(
        \add_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [1]), .IN2(\fadd_0_0_0_0_0/resultbeforeround [1]), .Q(
        \add_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [2]) );
  XOR2X1 U6965 ( .IN1(
        \add_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [1]), .IN2(\fadd_0_0_0_0_0/resultbeforeround [1]), .Q(
        \fadd_0_0_0_0_0/resultrounded [1]) );
  AND2X1 U6966 ( .IN1(\fadd_0_0_0_0_0/round ), .IN2(
        \fadd_0_0_0_0_0/resultbeforeround [0]), .Q(
        \add_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [1]) );
  XOR2X1 U6967 ( .IN1(\fadd_0_0_0_0_0/round ), .IN2(
        \fadd_0_0_0_0_0/resultbeforeround [0]), .Q(
        \fadd_0_0_0_0_0/resultrounded [0]) );
  AND2X1 U6968 ( .IN1(n14224), .IN2(\fadd_0_0_0_0_0/add_859/carry [5]), .Q(
        \fadd_0_0_0_0_0/add_859/carry [6]) );
  XOR2X1 U6969 ( .IN1(n14224), .IN2(\fadd_0_0_0_0_0/add_859/carry [5]), .Q(
        \fadd_0_0_0_0_0/exponentresultfar1 [5]) );
  AND2X1 U6970 ( .IN1(\fadd_0_0_0_0_0/expoperationsel[0] ), .IN2(
        \fadd_0_0_0_0_0/exponentresultfar0_d2 [0]), .Q(
        \fadd_0_0_0_0_0/add_859/carry [1]) );
  XOR2X1 U6971 ( .IN1(\fadd_0_0_0_0_0/expoperationsel[0] ), .IN2(
        \fadd_0_0_0_0_0/exponentresultfar0_d2 [0]), .Q(
        \fadd_0_0_0_0_0/exponentresultfar1 [0]) );
  XNOR2X1 U6972 ( .IN1(\fadd_0_0_0_0_4/newx_d1 [8]), .IN2(
        \fadd_0_0_0_0_4/sub_784/carry [4]), .Q(
        \fadd_0_0_0_0_4/exponentresultclose [4]) );
  OR2X1 U6973 ( .IN1(\fadd_0_0_0_0_4/sub_784/carry [3]), .IN2(
        \fadd_0_0_0_0_4/newx_d1 [7]), .Q(\fadd_0_0_0_0_4/sub_784/carry [4]) );
  XNOR2X1 U6974 ( .IN1(\fadd_0_0_0_0_4/newx_d1 [7]), .IN2(
        \fadd_0_0_0_0_4/sub_784/carry [3]), .Q(
        \fadd_0_0_0_0_4/exponentresultclose [3]) );
  OR2X1 U6975 ( .IN1(n14585), .IN2(\fadd_0_0_0_0_4/newx_d1 [4]), .Q(
        \fadd_0_0_0_0_4/sub_784/carry [1]) );
  XNOR2X1 U6976 ( .IN1(\fadd_0_0_0_0_4/newx_d1 [4]), .IN2(n14585), .Q(
        \fadd_0_0_0_0_4/exponentresultclose [0]) );
  XOR2X1 U6977 ( .IN1(
        \add_1_root_fmul_0_0_0_0_0/roundingadder/add_57/carry [10]), .IN2(
        \fmul_0_0_0_0_0/roundingadder/x_1_d1 [10]), .Q(
        \fmul_0_0_0_0_0/expsigpostround [10]) );
  AND2X1 U6978 ( .IN1(
        \add_1_root_fmul_0_0_0_0_0/roundingadder/add_57/carry [9]), .IN2(
        \fmul_0_0_0_0_0/roundingadder/x_1_d1 [9]), .Q(
        \add_1_root_fmul_0_0_0_0_0/roundingadder/add_57/carry [10]) );
  XOR2X1 U6979 ( .IN1(
        \add_1_root_fmul_0_0_0_0_0/roundingadder/add_57/carry [9]), .IN2(
        \fmul_0_0_0_0_0/roundingadder/x_1_d1 [9]), .Q(
        \fmul_0_0_0_0_0/expsigpostround [9]) );
  AND2X1 U6980 ( .IN1(\fmul_0_0_0_0_0/roundingadder/x_1_d1 [8]), .IN2(
        \add_1_root_fmul_0_0_0_0_0/roundingadder/add_57/carry [8]), .Q(
        \add_1_root_fmul_0_0_0_0_0/roundingadder/add_57/carry [9]) );
  XOR2X1 U6981 ( .IN1(
        \add_1_root_fmul_0_0_0_0_0/roundingadder/add_57/carry [8]), .IN2(
        \fmul_0_0_0_0_0/roundingadder/x_1_d1 [8]), .Q(\U565/DATA2_8 ) );
  AND2X1 U6982 ( .IN1(\fmul_0_0_0_0_0/roundingadder/x_1_d1 [7]), .IN2(
        \add_1_root_fmul_0_0_0_0_0/roundingadder/add_57/carry [7]), .Q(
        \add_1_root_fmul_0_0_0_0_0/roundingadder/add_57/carry [8]) );
  XOR2X1 U6983 ( .IN1(
        \add_1_root_fmul_0_0_0_0_0/roundingadder/add_57/carry [7]), .IN2(
        \fmul_0_0_0_0_0/roundingadder/x_1_d1 [7]), .Q(\U565/DATA2_7 ) );
  AND2X1 U6984 ( .IN1(\fmul_0_0_0_0_0/roundingadder/x_1_d1 [6]), .IN2(
        \add_1_root_fmul_0_0_0_0_0/roundingadder/add_57/carry [6]), .Q(
        \add_1_root_fmul_0_0_0_0_0/roundingadder/add_57/carry [7]) );
  XOR2X1 U6985 ( .IN1(
        \add_1_root_fmul_0_0_0_0_0/roundingadder/add_57/carry [6]), .IN2(
        \fmul_0_0_0_0_0/roundingadder/x_1_d1 [6]), .Q(\U565/DATA2_6 ) );
  AND2X1 U6986 ( .IN1(\fmul_0_0_0_0_0/roundingadder/x_1_d1 [5]), .IN2(
        \add_1_root_fmul_0_0_0_0_0/roundingadder/add_57/carry [5]), .Q(
        \add_1_root_fmul_0_0_0_0_0/roundingadder/add_57/carry [6]) );
  XOR2X1 U6987 ( .IN1(
        \add_1_root_fmul_0_0_0_0_0/roundingadder/add_57/carry [5]), .IN2(
        \fmul_0_0_0_0_0/roundingadder/x_1_d1 [5]), .Q(\U565/DATA2_5 ) );
  AND2X1 U6988 ( .IN1(\fmul_0_0_0_0_0/roundingadder/x_1_d1 [4]), .IN2(
        \add_1_root_fmul_0_0_0_0_0/roundingadder/add_57/carry [4]), .Q(
        \add_1_root_fmul_0_0_0_0_0/roundingadder/add_57/carry [5]) );
  XOR2X1 U6989 ( .IN1(
        \add_1_root_fmul_0_0_0_0_0/roundingadder/add_57/carry [4]), .IN2(
        \fmul_0_0_0_0_0/roundingadder/x_1_d1 [4]), .Q(\U565/DATA2_4 ) );
  AND2X1 U6990 ( .IN1(\fmul_0_0_0_0_0/roundingadder/x_1_d1 [3]), .IN2(
        \add_1_root_fmul_0_0_0_0_0/roundingadder/add_57/carry [3]), .Q(
        \add_1_root_fmul_0_0_0_0_0/roundingadder/add_57/carry [4]) );
  XOR2X1 U6991 ( .IN1(
        \add_1_root_fmul_0_0_0_0_0/roundingadder/add_57/carry [3]), .IN2(
        \fmul_0_0_0_0_0/roundingadder/x_1_d1 [3]), .Q(\U565/DATA2_3 ) );
  AND2X1 U6992 ( .IN1(\fmul_0_0_0_0_0/roundingadder/x_1_d1 [2]), .IN2(
        \add_1_root_fmul_0_0_0_0_0/roundingadder/add_57/carry [2]), .Q(
        \add_1_root_fmul_0_0_0_0_0/roundingadder/add_57/carry [3]) );
  XOR2X1 U6993 ( .IN1(
        \add_1_root_fmul_0_0_0_0_0/roundingadder/add_57/carry [2]), .IN2(
        \fmul_0_0_0_0_0/roundingadder/x_1_d1 [2]), .Q(\U565/DATA2_2 ) );
  AND2X1 U6994 ( .IN1(\fmul_0_0_0_0_0/roundingadder/x_1_d1 [1]), .IN2(
        \add_1_root_fmul_0_0_0_0_0/roundingadder/add_57/carry [1]), .Q(
        \add_1_root_fmul_0_0_0_0_0/roundingadder/add_57/carry [2]) );
  XOR2X1 U6995 ( .IN1(
        \add_1_root_fmul_0_0_0_0_0/roundingadder/add_57/carry [1]), .IN2(
        \fmul_0_0_0_0_0/roundingadder/x_1_d1 [1]), .Q(\U565/DATA2_1 ) );
  AND2X1 U6996 ( .IN1(\fmul_0_0_0_0_0/roundingadder/x_1_d1 [0]), .IN2(
        \fmul_0_0_0_0_0/roundingadder/n151_o[0] ), .Q(
        \add_1_root_fmul_0_0_0_0_0/roundingadder/add_57/carry [1]) );
  XOR2X1 U6997 ( .IN1(\fmul_0_0_0_0_0/roundingadder/n151_o[0] ), .IN2(
        \fmul_0_0_0_0_0/roundingadder/x_1_d1 [0]), .Q(\U565/DATA2_0 ) );
  XOR2X1 U6998 ( .IN1(
        \add_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [10]), .IN2(\fadd_0_0_0_0_4/resultbeforeround [10]), .Q(
        \fadd_0_0_0_0_4/resultrounded [10]) );
  XOR2X1 U6999 ( .IN1(n14228), .IN2(\fadd_0_0_0_0_4/add_859/carry [6]), .Q(
        \fadd_0_0_0_0_4/exponentresultfar1 [6]) );
  AND2X1 U7000 ( .IN1(
        \add_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [9]), .IN2(\fadd_0_0_0_0_4/resultbeforeround [9]), .Q(
        \add_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [10]) );
  AND2X1 U7001 ( .IN1(
        \add_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [8]), .IN2(\fadd_0_0_0_0_4/resultbeforeround [8]), .Q(
        \add_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [9]) );
  XOR2X1 U7002 ( .IN1(
        \add_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [8]), .IN2(\fadd_0_0_0_0_4/resultbeforeround [8]), .Q(
        \fadd_0_0_0_0_4/resultrounded [8]) );
  AND2X1 U7003 ( .IN1(
        \add_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [7]), .IN2(\fadd_0_0_0_0_4/resultbeforeround [7]), .Q(
        \add_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [8]) );
  XOR2X1 U7004 ( .IN1(
        \add_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [7]), .IN2(\fadd_0_0_0_0_4/resultbeforeround [7]), .Q(
        \fadd_0_0_0_0_4/resultrounded [7]) );
  AND2X1 U7005 ( .IN1(
        \add_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [6]), .IN2(\fadd_0_0_0_0_4/resultbeforeround [6]), .Q(
        \add_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [7]) );
  XOR2X1 U7006 ( .IN1(
        \add_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [6]), .IN2(\fadd_0_0_0_0_4/resultbeforeround [6]), .Q(
        \fadd_0_0_0_0_4/resultrounded [6]) );
  AND2X1 U7007 ( .IN1(
        \add_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [5]), .IN2(\fadd_0_0_0_0_4/resultbeforeround [5]), .Q(
        \add_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [6]) );
  XOR2X1 U7008 ( .IN1(
        \add_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [5]), .IN2(\fadd_0_0_0_0_4/resultbeforeround [5]), .Q(
        \fadd_0_0_0_0_4/resultrounded [5]) );
  AND2X1 U7009 ( .IN1(
        \add_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [4]), .IN2(\fadd_0_0_0_0_4/resultbeforeround [4]), .Q(
        \add_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [5]) );
  XOR2X1 U7010 ( .IN1(
        \add_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [4]), .IN2(\fadd_0_0_0_0_4/resultbeforeround [4]), .Q(
        \fadd_0_0_0_0_4/resultrounded [4]) );
  AND2X1 U7011 ( .IN1(
        \add_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [3]), .IN2(\fadd_0_0_0_0_4/resultbeforeround [3]), .Q(
        \add_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [4]) );
  XOR2X1 U7012 ( .IN1(
        \add_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [3]), .IN2(\fadd_0_0_0_0_4/resultbeforeround [3]), .Q(
        \fadd_0_0_0_0_4/resultrounded [3]) );
  AND2X1 U7013 ( .IN1(
        \add_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [2]), .IN2(\fadd_0_0_0_0_4/resultbeforeround [2]), .Q(
        \add_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [3]) );
  XOR2X1 U7014 ( .IN1(
        \add_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [2]), .IN2(\fadd_0_0_0_0_4/resultbeforeround [2]), .Q(
        \fadd_0_0_0_0_4/resultrounded [2]) );
  AND2X1 U7015 ( .IN1(
        \add_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [1]), .IN2(\fadd_0_0_0_0_4/resultbeforeround [1]), .Q(
        \add_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [2]) );
  XOR2X1 U7016 ( .IN1(
        \add_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [1]), .IN2(\fadd_0_0_0_0_4/resultbeforeround [1]), .Q(
        \fadd_0_0_0_0_4/resultrounded [1]) );
  AND2X1 U7017 ( .IN1(\fadd_0_0_0_0_4/round ), .IN2(
        \fadd_0_0_0_0_4/resultbeforeround [0]), .Q(
        \add_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [1]) );
  XOR2X1 U7018 ( .IN1(\fadd_0_0_0_0_4/round ), .IN2(
        \fadd_0_0_0_0_4/resultbeforeround [0]), .Q(
        \fadd_0_0_0_0_4/resultrounded [0]) );
  AND2X1 U7019 ( .IN1(n14228), .IN2(\fadd_0_0_0_0_4/add_859/carry [5]), .Q(
        \fadd_0_0_0_0_4/add_859/carry [6]) );
  XOR2X1 U7020 ( .IN1(n14228), .IN2(\fadd_0_0_0_0_4/add_859/carry [5]), .Q(
        \fadd_0_0_0_0_4/exponentresultfar1 [5]) );
  AND2X1 U7021 ( .IN1(\fadd_0_0_0_0_4/expoperationsel[0] ), .IN2(
        \fadd_0_0_0_0_4/exponentresultfar0_d2 [0]), .Q(
        \fadd_0_0_0_0_4/add_859/carry [1]) );
  XOR2X1 U7022 ( .IN1(\fadd_0_0_0_0_4/expoperationsel[0] ), .IN2(
        \fadd_0_0_0_0_4/exponentresultfar0_d2 [0]), .Q(
        \fadd_0_0_0_0_4/exponentresultfar1 [0]) );
  XNOR2X1 U7023 ( .IN1(\fadd_0_0_0_0_6/newx_d1 [8]), .IN2(
        \fadd_0_0_0_0_6/sub_784/carry [4]), .Q(
        \fadd_0_0_0_0_6/exponentresultclose [4]) );
  OR2X1 U7024 ( .IN1(\fadd_0_0_0_0_6/sub_784/carry [3]), .IN2(
        \fadd_0_0_0_0_6/newx_d1 [7]), .Q(\fadd_0_0_0_0_6/sub_784/carry [4]) );
  XNOR2X1 U7025 ( .IN1(\fadd_0_0_0_0_6/newx_d1 [7]), .IN2(
        \fadd_0_0_0_0_6/sub_784/carry [3]), .Q(
        \fadd_0_0_0_0_6/exponentresultclose [3]) );
  OR2X1 U7026 ( .IN1(n14607), .IN2(\fadd_0_0_0_0_6/newx_d1 [4]), .Q(
        \fadd_0_0_0_0_6/sub_784/carry [1]) );
  XNOR2X1 U7027 ( .IN1(\fadd_0_0_0_0_6/newx_d1 [4]), .IN2(n14607), .Q(
        \fadd_0_0_0_0_6/exponentresultclose [0]) );
  XOR2X1 U7028 ( .IN1(
        \add_1_root_fmul_0_0_0_0_4/roundingadder/add_57/carry [10]), .IN2(
        \fmul_0_0_0_0_4/roundingadder/x_1_d1 [10]), .Q(
        \fmul_0_0_0_0_4/expsigpostround [10]) );
  AND2X1 U7029 ( .IN1(
        \add_1_root_fmul_0_0_0_0_4/roundingadder/add_57/carry [9]), .IN2(
        \fmul_0_0_0_0_4/roundingadder/x_1_d1 [9]), .Q(
        \add_1_root_fmul_0_0_0_0_4/roundingadder/add_57/carry [10]) );
  XOR2X1 U7030 ( .IN1(
        \add_1_root_fmul_0_0_0_0_4/roundingadder/add_57/carry [9]), .IN2(
        \fmul_0_0_0_0_4/roundingadder/x_1_d1 [9]), .Q(
        \fmul_0_0_0_0_4/expsigpostround [9]) );
  AND2X1 U7031 ( .IN1(\fmul_0_0_0_0_4/roundingadder/x_1_d1 [8]), .IN2(
        \add_1_root_fmul_0_0_0_0_4/roundingadder/add_57/carry [8]), .Q(
        \add_1_root_fmul_0_0_0_0_4/roundingadder/add_57/carry [9]) );
  XOR2X1 U7032 ( .IN1(
        \add_1_root_fmul_0_0_0_0_4/roundingadder/add_57/carry [8]), .IN2(
        \fmul_0_0_0_0_4/roundingadder/x_1_d1 [8]), .Q(\U341/DATA2_8 ) );
  AND2X1 U7033 ( .IN1(\fmul_0_0_0_0_4/roundingadder/x_1_d1 [7]), .IN2(
        \add_1_root_fmul_0_0_0_0_4/roundingadder/add_57/carry [7]), .Q(
        \add_1_root_fmul_0_0_0_0_4/roundingadder/add_57/carry [8]) );
  XOR2X1 U7034 ( .IN1(
        \add_1_root_fmul_0_0_0_0_4/roundingadder/add_57/carry [7]), .IN2(
        \fmul_0_0_0_0_4/roundingadder/x_1_d1 [7]), .Q(\U341/DATA2_7 ) );
  AND2X1 U7035 ( .IN1(\fmul_0_0_0_0_4/roundingadder/x_1_d1 [6]), .IN2(
        \add_1_root_fmul_0_0_0_0_4/roundingadder/add_57/carry [6]), .Q(
        \add_1_root_fmul_0_0_0_0_4/roundingadder/add_57/carry [7]) );
  XOR2X1 U7036 ( .IN1(
        \add_1_root_fmul_0_0_0_0_4/roundingadder/add_57/carry [6]), .IN2(
        \fmul_0_0_0_0_4/roundingadder/x_1_d1 [6]), .Q(\U341/DATA2_6 ) );
  AND2X1 U7037 ( .IN1(\fmul_0_0_0_0_4/roundingadder/x_1_d1 [5]), .IN2(
        \add_1_root_fmul_0_0_0_0_4/roundingadder/add_57/carry [5]), .Q(
        \add_1_root_fmul_0_0_0_0_4/roundingadder/add_57/carry [6]) );
  XOR2X1 U7038 ( .IN1(
        \add_1_root_fmul_0_0_0_0_4/roundingadder/add_57/carry [5]), .IN2(
        \fmul_0_0_0_0_4/roundingadder/x_1_d1 [5]), .Q(\U341/DATA2_5 ) );
  AND2X1 U7039 ( .IN1(\fmul_0_0_0_0_4/roundingadder/x_1_d1 [4]), .IN2(
        \add_1_root_fmul_0_0_0_0_4/roundingadder/add_57/carry [4]), .Q(
        \add_1_root_fmul_0_0_0_0_4/roundingadder/add_57/carry [5]) );
  XOR2X1 U7040 ( .IN1(
        \add_1_root_fmul_0_0_0_0_4/roundingadder/add_57/carry [4]), .IN2(
        \fmul_0_0_0_0_4/roundingadder/x_1_d1 [4]), .Q(\U341/DATA2_4 ) );
  AND2X1 U7041 ( .IN1(\fmul_0_0_0_0_4/roundingadder/x_1_d1 [3]), .IN2(
        \add_1_root_fmul_0_0_0_0_4/roundingadder/add_57/carry [3]), .Q(
        \add_1_root_fmul_0_0_0_0_4/roundingadder/add_57/carry [4]) );
  XOR2X1 U7042 ( .IN1(
        \add_1_root_fmul_0_0_0_0_4/roundingadder/add_57/carry [3]), .IN2(
        \fmul_0_0_0_0_4/roundingadder/x_1_d1 [3]), .Q(\U341/DATA2_3 ) );
  AND2X1 U7043 ( .IN1(\fmul_0_0_0_0_4/roundingadder/x_1_d1 [2]), .IN2(
        \add_1_root_fmul_0_0_0_0_4/roundingadder/add_57/carry [2]), .Q(
        \add_1_root_fmul_0_0_0_0_4/roundingadder/add_57/carry [3]) );
  XOR2X1 U7044 ( .IN1(
        \add_1_root_fmul_0_0_0_0_4/roundingadder/add_57/carry [2]), .IN2(
        \fmul_0_0_0_0_4/roundingadder/x_1_d1 [2]), .Q(\U341/DATA2_2 ) );
  AND2X1 U7045 ( .IN1(\fmul_0_0_0_0_4/roundingadder/x_1_d1 [1]), .IN2(
        \add_1_root_fmul_0_0_0_0_4/roundingadder/add_57/carry [1]), .Q(
        \add_1_root_fmul_0_0_0_0_4/roundingadder/add_57/carry [2]) );
  XOR2X1 U7046 ( .IN1(
        \add_1_root_fmul_0_0_0_0_4/roundingadder/add_57/carry [1]), .IN2(
        \fmul_0_0_0_0_4/roundingadder/x_1_d1 [1]), .Q(\U341/DATA2_1 ) );
  AND2X1 U7047 ( .IN1(\fmul_0_0_0_0_4/roundingadder/n151_o[0] ), .IN2(
        \fmul_0_0_0_0_4/roundingadder/x_1_d1 [0]), .Q(
        \add_1_root_fmul_0_0_0_0_4/roundingadder/add_57/carry [1]) );
  XOR2X1 U7048 ( .IN1(\fmul_0_0_0_0_4/roundingadder/n151_o[0] ), .IN2(
        \fmul_0_0_0_0_4/roundingadder/x_1_d1 [0]), .Q(n13466) );
  XOR2X1 U7049 ( .IN1(
        \add_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [10]), .IN2(\fadd_0_0_0_0_6/resultbeforeround [10]), .Q(
        \fadd_0_0_0_0_6/resultrounded [10]) );
  XOR2X1 U7050 ( .IN1(\fadd_0_0_0_0_6/add_859/B[1] ), .IN2(
        \fadd_0_0_0_0_6/add_859/carry [6]), .Q(
        \fadd_0_0_0_0_6/exponentresultfar1 [6]) );
  AND2X1 U7051 ( .IN1(
        \add_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [9]), .IN2(\fadd_0_0_0_0_6/resultbeforeround [9]), .Q(
        \add_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [10]) );
  XOR2X1 U7052 ( .IN1(
        \add_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [9]), .IN2(\fadd_0_0_0_0_6/resultbeforeround [9]), .Q(
        \fadd_0_0_0_0_6/resultrounded [9]) );
  AND2X1 U7053 ( .IN1(
        \add_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [8]), .IN2(\fadd_0_0_0_0_6/resultbeforeround [8]), .Q(
        \add_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [9]) );
  XOR2X1 U7054 ( .IN1(
        \add_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [8]), .IN2(\fadd_0_0_0_0_6/resultbeforeround [8]), .Q(
        \fadd_0_0_0_0_6/resultrounded [8]) );
  AND2X1 U7055 ( .IN1(
        \add_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [7]), .IN2(\fadd_0_0_0_0_6/resultbeforeround [7]), .Q(
        \add_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [8]) );
  XOR2X1 U7056 ( .IN1(
        \add_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [7]), .IN2(\fadd_0_0_0_0_6/resultbeforeround [7]), .Q(
        \fadd_0_0_0_0_6/resultrounded [7]) );
  AND2X1 U7057 ( .IN1(
        \add_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [6]), .IN2(\fadd_0_0_0_0_6/resultbeforeround [6]), .Q(
        \add_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [7]) );
  XOR2X1 U7058 ( .IN1(
        \add_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [6]), .IN2(\fadd_0_0_0_0_6/resultbeforeround [6]), .Q(
        \fadd_0_0_0_0_6/resultrounded [6]) );
  AND2X1 U7059 ( .IN1(
        \add_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [5]), .IN2(\fadd_0_0_0_0_6/resultbeforeround [5]), .Q(
        \add_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [6]) );
  XOR2X1 U7060 ( .IN1(
        \add_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [5]), .IN2(\fadd_0_0_0_0_6/resultbeforeround [5]), .Q(
        \fadd_0_0_0_0_6/resultrounded [5]) );
  AND2X1 U7061 ( .IN1(
        \add_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [4]), .IN2(\fadd_0_0_0_0_6/resultbeforeround [4]), .Q(
        \add_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [5]) );
  XOR2X1 U7062 ( .IN1(
        \add_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [4]), .IN2(\fadd_0_0_0_0_6/resultbeforeround [4]), .Q(
        \fadd_0_0_0_0_6/resultrounded [4]) );
  AND2X1 U7063 ( .IN1(
        \add_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [3]), .IN2(\fadd_0_0_0_0_6/resultbeforeround [3]), .Q(
        \add_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [4]) );
  XOR2X1 U7064 ( .IN1(
        \add_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [3]), .IN2(\fadd_0_0_0_0_6/resultbeforeround [3]), .Q(
        \fadd_0_0_0_0_6/resultrounded [3]) );
  AND2X1 U7065 ( .IN1(
        \add_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [2]), .IN2(\fadd_0_0_0_0_6/resultbeforeround [2]), .Q(
        \add_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [3]) );
  XOR2X1 U7066 ( .IN1(
        \add_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [2]), .IN2(\fadd_0_0_0_0_6/resultbeforeround [2]), .Q(
        \fadd_0_0_0_0_6/resultrounded [2]) );
  AND2X1 U7067 ( .IN1(
        \add_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [1]), .IN2(\fadd_0_0_0_0_6/resultbeforeround [1]), .Q(
        \add_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [2]) );
  XOR2X1 U7068 ( .IN1(
        \add_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [1]), .IN2(\fadd_0_0_0_0_6/resultbeforeround [1]), .Q(
        \fadd_0_0_0_0_6/resultrounded [1]) );
  AND2X1 U7069 ( .IN1(\fadd_0_0_0_0_6/round ), .IN2(
        \fadd_0_0_0_0_6/resultbeforeround [0]), .Q(
        \add_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [1]) );
  XOR2X1 U7070 ( .IN1(\fadd_0_0_0_0_6/round ), .IN2(
        \fadd_0_0_0_0_6/resultbeforeround [0]), .Q(
        \fadd_0_0_0_0_6/resultrounded [0]) );
  AND2X1 U7071 ( .IN1(\fadd_0_0_0_0_6/add_859/B[1] ), .IN2(
        \fadd_0_0_0_0_6/add_859/carry [5]), .Q(
        \fadd_0_0_0_0_6/add_859/carry [6]) );
  XOR2X1 U7072 ( .IN1(\fadd_0_0_0_0_6/add_859/B[1] ), .IN2(
        \fadd_0_0_0_0_6/add_859/carry [5]), .Q(
        \fadd_0_0_0_0_6/exponentresultfar1 [5]) );
  AND2X1 U7073 ( .IN1(\fadd_0_0_0_0_6/expoperationsel[0] ), .IN2(
        \fadd_0_0_0_0_6/exponentresultfar0_d2 [0]), .Q(
        \fadd_0_0_0_0_6/add_859/carry [1]) );
  XOR2X1 U7074 ( .IN1(\fadd_0_0_0_0_6/expoperationsel[0] ), .IN2(
        \fadd_0_0_0_0_6/exponentresultfar0_d2 [0]), .Q(
        \fadd_0_0_0_0_6/exponentresultfar1 [0]) );
  XNOR2X1 U7075 ( .IN1(\fadd_0_0_0_0_7/newx_d1 [8]), .IN2(
        \fadd_0_0_0_0_7/sub_784/carry [4]), .Q(
        \fadd_0_0_0_0_7/exponentresultclose [4]) );
  OR2X1 U7076 ( .IN1(\fadd_0_0_0_0_7/sub_784/carry [3]), .IN2(
        \fadd_0_0_0_0_7/newx_d1 [7]), .Q(\fadd_0_0_0_0_7/sub_784/carry [4]) );
  XNOR2X1 U7077 ( .IN1(\fadd_0_0_0_0_7/newx_d1 [7]), .IN2(
        \fadd_0_0_0_0_7/sub_784/carry [3]), .Q(
        \fadd_0_0_0_0_7/exponentresultclose [3]) );
  OR2X1 U7078 ( .IN1(n14618), .IN2(\fadd_0_0_0_0_7/newx_d1 [4]), .Q(
        \fadd_0_0_0_0_7/sub_784/carry [1]) );
  XNOR2X1 U7079 ( .IN1(\fadd_0_0_0_0_7/newx_d1 [4]), .IN2(n14618), .Q(
        \fadd_0_0_0_0_7/exponentresultclose [0]) );
  XOR2X1 U7080 ( .IN1(
        \add_1_root_fmul_0_0_0_0_6/roundingadder/add_57/carry [10]), .IN2(
        \fmul_0_0_0_0_6/roundingadder/x_1_d1 [10]), .Q(
        \fmul_0_0_0_0_6/expsigpostround [10]) );
  AND2X1 U7081 ( .IN1(
        \add_1_root_fmul_0_0_0_0_6/roundingadder/add_57/carry [9]), .IN2(
        \fmul_0_0_0_0_6/roundingadder/x_1_d1 [9]), .Q(
        \add_1_root_fmul_0_0_0_0_6/roundingadder/add_57/carry [10]) );
  XOR2X1 U7082 ( .IN1(
        \add_1_root_fmul_0_0_0_0_6/roundingadder/add_57/carry [9]), .IN2(
        \fmul_0_0_0_0_6/roundingadder/x_1_d1 [9]), .Q(
        \fmul_0_0_0_0_6/expsigpostround [9]) );
  AND2X1 U7083 ( .IN1(\fmul_0_0_0_0_6/roundingadder/x_1_d1 [8]), .IN2(
        \add_1_root_fmul_0_0_0_0_6/roundingadder/add_57/carry [8]), .Q(
        \add_1_root_fmul_0_0_0_0_6/roundingadder/add_57/carry [9]) );
  XOR2X1 U7084 ( .IN1(
        \add_1_root_fmul_0_0_0_0_6/roundingadder/add_57/carry [8]), .IN2(
        \fmul_0_0_0_0_6/roundingadder/x_1_d1 [8]), .Q(\U229/DATA2_8 ) );
  AND2X1 U7085 ( .IN1(\fmul_0_0_0_0_6/roundingadder/x_1_d1 [7]), .IN2(
        \add_1_root_fmul_0_0_0_0_6/roundingadder/add_57/carry [7]), .Q(
        \add_1_root_fmul_0_0_0_0_6/roundingadder/add_57/carry [8]) );
  XOR2X1 U7086 ( .IN1(
        \add_1_root_fmul_0_0_0_0_6/roundingadder/add_57/carry [7]), .IN2(
        \fmul_0_0_0_0_6/roundingadder/x_1_d1 [7]), .Q(\U229/DATA2_7 ) );
  AND2X1 U7087 ( .IN1(\fmul_0_0_0_0_6/roundingadder/x_1_d1 [6]), .IN2(
        \add_1_root_fmul_0_0_0_0_6/roundingadder/add_57/carry [6]), .Q(
        \add_1_root_fmul_0_0_0_0_6/roundingadder/add_57/carry [7]) );
  XOR2X1 U7088 ( .IN1(
        \add_1_root_fmul_0_0_0_0_6/roundingadder/add_57/carry [6]), .IN2(
        \fmul_0_0_0_0_6/roundingadder/x_1_d1 [6]), .Q(\U229/DATA2_6 ) );
  AND2X1 U7089 ( .IN1(
        \add_1_root_fmul_0_0_0_0_6/roundingadder/add_57/carry [5]), .IN2(
        \fmul_0_0_0_0_6/roundingadder/x_1_d1 [5]), .Q(
        \add_1_root_fmul_0_0_0_0_6/roundingadder/add_57/carry [6]) );
  XOR2X1 U7090 ( .IN1(
        \add_1_root_fmul_0_0_0_0_6/roundingadder/add_57/carry [5]), .IN2(
        \fmul_0_0_0_0_6/roundingadder/x_1_d1 [5]), .Q(n13459) );
  AND2X1 U7091 ( .IN1(
        \add_1_root_fmul_0_0_0_0_6/roundingadder/add_57/carry [4]), .IN2(
        \fmul_0_0_0_0_6/roundingadder/x_1_d1 [4]), .Q(
        \add_1_root_fmul_0_0_0_0_6/roundingadder/add_57/carry [5]) );
  XOR2X1 U7092 ( .IN1(
        \add_1_root_fmul_0_0_0_0_6/roundingadder/add_57/carry [4]), .IN2(
        \fmul_0_0_0_0_6/roundingadder/x_1_d1 [4]), .Q(n13460) );
  AND2X1 U7093 ( .IN1(
        \add_1_root_fmul_0_0_0_0_6/roundingadder/add_57/carry [3]), .IN2(
        \fmul_0_0_0_0_6/roundingadder/x_1_d1 [3]), .Q(
        \add_1_root_fmul_0_0_0_0_6/roundingadder/add_57/carry [4]) );
  XOR2X1 U7094 ( .IN1(
        \add_1_root_fmul_0_0_0_0_6/roundingadder/add_57/carry [3]), .IN2(
        \fmul_0_0_0_0_6/roundingadder/x_1_d1 [3]), .Q(n13461) );
  AND2X1 U7095 ( .IN1(
        \add_1_root_fmul_0_0_0_0_6/roundingadder/add_57/carry [2]), .IN2(
        \fmul_0_0_0_0_6/roundingadder/x_1_d1 [2]), .Q(
        \add_1_root_fmul_0_0_0_0_6/roundingadder/add_57/carry [3]) );
  XOR2X1 U7096 ( .IN1(
        \add_1_root_fmul_0_0_0_0_6/roundingadder/add_57/carry [2]), .IN2(
        \fmul_0_0_0_0_6/roundingadder/x_1_d1 [2]), .Q(n13462) );
  AND2X1 U7097 ( .IN1(
        \add_1_root_fmul_0_0_0_0_6/roundingadder/add_57/carry [1]), .IN2(
        \fmul_0_0_0_0_6/roundingadder/x_1_d1 [1]), .Q(
        \add_1_root_fmul_0_0_0_0_6/roundingadder/add_57/carry [2]) );
  XOR2X1 U7098 ( .IN1(
        \add_1_root_fmul_0_0_0_0_6/roundingadder/add_57/carry [1]), .IN2(
        \fmul_0_0_0_0_6/roundingadder/x_1_d1 [1]), .Q(n13463) );
  XOR2X1 U7099 ( .IN1(
        \add_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [10]), .IN2(\fadd_0_0_0_0_7/resultbeforeround [10]), .Q(
        \fadd_0_0_0_0_7/resultrounded [10]) );
  XOR2X1 U7100 ( .IN1(n14231), .IN2(\fadd_0_0_0_0_7/add_859/carry [6]), .Q(
        \fadd_0_0_0_0_7/exponentresultfar1 [6]) );
  AND2X1 U7101 ( .IN1(
        \add_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [9]), .IN2(\fadd_0_0_0_0_7/resultbeforeround [9]), .Q(
        \add_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [10]) );
  XOR2X1 U7102 ( .IN1(
        \add_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [9]), .IN2(\fadd_0_0_0_0_7/resultbeforeround [9]), .Q(
        \fadd_0_0_0_0_7/resultrounded [9]) );
  AND2X1 U7103 ( .IN1(
        \add_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [8]), .IN2(\fadd_0_0_0_0_7/resultbeforeround [8]), .Q(
        \add_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [9]) );
  XOR2X1 U7104 ( .IN1(
        \add_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [8]), .IN2(\fadd_0_0_0_0_7/resultbeforeround [8]), .Q(
        \fadd_0_0_0_0_7/resultrounded [8]) );
  AND2X1 U7105 ( .IN1(
        \add_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [7]), .IN2(\fadd_0_0_0_0_7/resultbeforeround [7]), .Q(
        \add_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [8]) );
  XOR2X1 U7106 ( .IN1(
        \add_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [7]), .IN2(\fadd_0_0_0_0_7/resultbeforeround [7]), .Q(
        \fadd_0_0_0_0_7/resultrounded [7]) );
  AND2X1 U7107 ( .IN1(
        \add_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [6]), .IN2(\fadd_0_0_0_0_7/resultbeforeround [6]), .Q(
        \add_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [7]) );
  XOR2X1 U7108 ( .IN1(
        \add_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [6]), .IN2(\fadd_0_0_0_0_7/resultbeforeround [6]), .Q(
        \fadd_0_0_0_0_7/resultrounded [6]) );
  AND2X1 U7109 ( .IN1(
        \add_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [5]), .IN2(\fadd_0_0_0_0_7/resultbeforeround [5]), .Q(
        \add_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [6]) );
  XOR2X1 U7110 ( .IN1(
        \add_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [5]), .IN2(\fadd_0_0_0_0_7/resultbeforeround [5]), .Q(
        \fadd_0_0_0_0_7/resultrounded [5]) );
  AND2X1 U7111 ( .IN1(
        \add_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [4]), .IN2(\fadd_0_0_0_0_7/resultbeforeround [4]), .Q(
        \add_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [5]) );
  XOR2X1 U7112 ( .IN1(
        \add_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [4]), .IN2(\fadd_0_0_0_0_7/resultbeforeround [4]), .Q(
        \fadd_0_0_0_0_7/resultrounded [4]) );
  AND2X1 U7113 ( .IN1(
        \add_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [3]), .IN2(\fadd_0_0_0_0_7/resultbeforeround [3]), .Q(
        \add_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [4]) );
  XOR2X1 U7114 ( .IN1(
        \add_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [3]), .IN2(\fadd_0_0_0_0_7/resultbeforeround [3]), .Q(
        \fadd_0_0_0_0_7/resultrounded [3]) );
  AND2X1 U7115 ( .IN1(
        \add_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [2]), .IN2(\fadd_0_0_0_0_7/resultbeforeround [2]), .Q(
        \add_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [3]) );
  XOR2X1 U7116 ( .IN1(
        \add_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [2]), .IN2(\fadd_0_0_0_0_7/resultbeforeround [2]), .Q(
        \fadd_0_0_0_0_7/resultrounded [2]) );
  AND2X1 U7117 ( .IN1(
        \add_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [1]), .IN2(\fadd_0_0_0_0_7/resultbeforeround [1]), .Q(
        \add_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [2]) );
  XOR2X1 U7118 ( .IN1(
        \add_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [1]), .IN2(\fadd_0_0_0_0_7/resultbeforeround [1]), .Q(
        \fadd_0_0_0_0_7/resultrounded [1]) );
  AND2X1 U7119 ( .IN1(n14231), .IN2(\fadd_0_0_0_0_7/add_859/carry [5]), .Q(
        \fadd_0_0_0_0_7/add_859/carry [6]) );
  XOR2X1 U7120 ( .IN1(n14231), .IN2(\fadd_0_0_0_0_7/add_859/carry [5]), .Q(
        \fadd_0_0_0_0_7/exponentresultfar1 [5]) );
  AND2X1 U7121 ( .IN1(\fadd_0_0_0_0_7/expoperationsel[0] ), .IN2(
        \fadd_0_0_0_0_7/exponentresultfar0_d2 [0]), .Q(
        \fadd_0_0_0_0_7/add_859/carry [1]) );
  XOR2X1 U7122 ( .IN1(\fadd_0_0_0_0_7/expoperationsel[0] ), .IN2(
        \fadd_0_0_0_0_7/exponentresultfar0_d2 [0]), .Q(
        \fadd_0_0_0_0_7/exponentresultfar1 [0]) );
  AND2X1 U7123 ( .IN1(\fmul_0_0_0_0_6/roundingadder/n151_o[0] ), .IN2(
        \fmul_0_0_0_0_6/roundingadder/x_1_d1 [0]), .Q(
        \add_1_root_fmul_0_0_0_0_6/roundingadder/add_57/carry [1]) );
  XOR2X1 U7124 ( .IN1(\fmul_0_0_0_0_6/roundingadder/n151_o[0] ), .IN2(
        \fmul_0_0_0_0_6/roundingadder/x_1_d1 [0]), .Q(n13464) );
  AND2X1 U7125 ( .IN1(\fadd_0_0_0_0_7/round ), .IN2(
        \fadd_0_0_0_0_7/resultbeforeround [0]), .Q(
        \add_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [1]) );
  XOR2X1 U7126 ( .IN1(\fadd_0_0_0_0_7/round ), .IN2(
        \fadd_0_0_0_0_7/resultbeforeround [0]), .Q(
        \fadd_0_0_0_0_7/resultrounded [0]) );
  XOR2X1 U7127 ( .IN1(
        \add_1_root_fmul_0_0_0_0_7/roundingadder/add_57/carry [10]), .IN2(
        \fmul_0_0_0_0_7/roundingadder/x_1_d1 [10]), .Q(
        \fmul_0_0_0_0_7/expsigpostround [10]) );
  AND2X1 U7128 ( .IN1(
        \add_1_root_fmul_0_0_0_0_7/roundingadder/add_57/carry [9]), .IN2(
        \fmul_0_0_0_0_7/roundingadder/x_1_d1 [9]), .Q(
        \add_1_root_fmul_0_0_0_0_7/roundingadder/add_57/carry [10]) );
  XOR2X1 U7129 ( .IN1(
        \add_1_root_fmul_0_0_0_0_7/roundingadder/add_57/carry [9]), .IN2(
        \fmul_0_0_0_0_7/roundingadder/x_1_d1 [9]), .Q(
        \fmul_0_0_0_0_7/expsigpostround [9]) );
  AND2X1 U7130 ( .IN1(\fmul_0_0_0_0_7/roundingadder/x_1_d1 [8]), .IN2(
        \add_1_root_fmul_0_0_0_0_7/roundingadder/add_57/carry [8]), .Q(
        \add_1_root_fmul_0_0_0_0_7/roundingadder/add_57/carry [9]) );
  XOR2X1 U7131 ( .IN1(
        \add_1_root_fmul_0_0_0_0_7/roundingadder/add_57/carry [8]), .IN2(
        \fmul_0_0_0_0_7/roundingadder/x_1_d1 [8]), .Q(\U173/DATA2_8 ) );
  AND2X1 U7132 ( .IN1(\fmul_0_0_0_0_7/roundingadder/x_1_d1 [7]), .IN2(
        \add_1_root_fmul_0_0_0_0_7/roundingadder/add_57/carry [7]), .Q(
        \add_1_root_fmul_0_0_0_0_7/roundingadder/add_57/carry [8]) );
  XOR2X1 U7133 ( .IN1(
        \add_1_root_fmul_0_0_0_0_7/roundingadder/add_57/carry [7]), .IN2(
        \fmul_0_0_0_0_7/roundingadder/x_1_d1 [7]), .Q(\U173/DATA2_7 ) );
  AND2X1 U7134 ( .IN1(\fmul_0_0_0_0_7/roundingadder/x_1_d1 [6]), .IN2(
        \add_1_root_fmul_0_0_0_0_7/roundingadder/add_57/carry [6]), .Q(
        \add_1_root_fmul_0_0_0_0_7/roundingadder/add_57/carry [7]) );
  XOR2X1 U7135 ( .IN1(
        \add_1_root_fmul_0_0_0_0_7/roundingadder/add_57/carry [6]), .IN2(
        \fmul_0_0_0_0_7/roundingadder/x_1_d1 [6]), .Q(\U173/DATA2_6 ) );
  AND2X1 U7136 ( .IN1(\fmul_0_0_0_0_7/roundingadder/x_1_d1 [5]), .IN2(
        \add_1_root_fmul_0_0_0_0_7/roundingadder/add_57/carry [5]), .Q(
        \add_1_root_fmul_0_0_0_0_7/roundingadder/add_57/carry [6]) );
  XOR2X1 U7137 ( .IN1(
        \add_1_root_fmul_0_0_0_0_7/roundingadder/add_57/carry [5]), .IN2(
        \fmul_0_0_0_0_7/roundingadder/x_1_d1 [5]), .Q(\U173/DATA2_5 ) );
  AND2X1 U7138 ( .IN1(\fmul_0_0_0_0_7/roundingadder/x_1_d1 [4]), .IN2(
        \add_1_root_fmul_0_0_0_0_7/roundingadder/add_57/carry [4]), .Q(
        \add_1_root_fmul_0_0_0_0_7/roundingadder/add_57/carry [5]) );
  XOR2X1 U7139 ( .IN1(
        \add_1_root_fmul_0_0_0_0_7/roundingadder/add_57/carry [4]), .IN2(
        \fmul_0_0_0_0_7/roundingadder/x_1_d1 [4]), .Q(\U173/DATA2_4 ) );
  AND2X1 U7140 ( .IN1(\fmul_0_0_0_0_7/roundingadder/x_1_d1 [3]), .IN2(
        \add_1_root_fmul_0_0_0_0_7/roundingadder/add_57/carry [3]), .Q(
        \add_1_root_fmul_0_0_0_0_7/roundingadder/add_57/carry [4]) );
  XOR2X1 U7141 ( .IN1(
        \add_1_root_fmul_0_0_0_0_7/roundingadder/add_57/carry [3]), .IN2(
        \fmul_0_0_0_0_7/roundingadder/x_1_d1 [3]), .Q(\U173/DATA2_3 ) );
  AND2X1 U7142 ( .IN1(\fmul_0_0_0_0_7/roundingadder/x_1_d1 [2]), .IN2(
        \add_1_root_fmul_0_0_0_0_7/roundingadder/add_57/carry [2]), .Q(
        \add_1_root_fmul_0_0_0_0_7/roundingadder/add_57/carry [3]) );
  XOR2X1 U7143 ( .IN1(
        \add_1_root_fmul_0_0_0_0_7/roundingadder/add_57/carry [2]), .IN2(
        \fmul_0_0_0_0_7/roundingadder/x_1_d1 [2]), .Q(\U173/DATA2_2 ) );
  AND2X1 U7144 ( .IN1(
        \add_1_root_fmul_0_0_0_0_7/roundingadder/add_57/carry [1]), .IN2(
        \fmul_0_0_0_0_7/roundingadder/x_1_d1 [1]), .Q(
        \add_1_root_fmul_0_0_0_0_7/roundingadder/add_57/carry [2]) );
  XOR2X1 U7145 ( .IN1(
        \add_1_root_fmul_0_0_0_0_7/roundingadder/add_57/carry [1]), .IN2(
        \fmul_0_0_0_0_7/roundingadder/x_1_d1 [1]), .Q(n13457) );
  AND2X1 U7146 ( .IN1(\fmul_0_0_0_0_7/roundingadder/n151_o[0] ), .IN2(
        \fmul_0_0_0_0_7/roundingadder/x_1_d1 [0]), .Q(
        \add_1_root_fmul_0_0_0_0_7/roundingadder/add_57/carry [1]) );
  XOR2X1 U7147 ( .IN1(\fmul_0_0_0_0_7/roundingadder/n151_o[0] ), .IN2(
        \fmul_0_0_0_0_7/roundingadder/x_1_d1 [0]), .Q(n13458) );
  XNOR2X1 U7148 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/A[5] ), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/carry [5]), .Q(
        \fmul_0_0_0_0_7/exppostnorm [5]) );
  OR2X1 U7149 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/carry [4]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/A[4] ), .Q(
        \add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/carry [5]) );
  XNOR2X1 U7150 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/A[4] ), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/carry [4]), .Q(
        \fmul_0_0_0_0_7/exppostnorm [4]) );
  AND2X1 U7151 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/carry [3]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/A[3] ), .Q(
        \add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/carry [4]) );
  XOR2X1 U7152 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/carry [3]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/A[3] ), .Q(
        \fmul_0_0_0_0_7/exppostnorm [3]) );
  AND2X1 U7153 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/carry [2]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/A[2] ), .Q(
        \add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/carry [3]) );
  XOR2X1 U7154 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/carry [2]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/A[2] ), .Q(
        \fmul_0_0_0_0_7/exppostnorm [2]) );
  AND2X1 U7155 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/B[0] ), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/A[0] ), .Q(
        \add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/carry [1]) );
  XOR2X1 U7156 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/B[0] ), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/A[0] ), .Q(
        \fmul_0_0_0_0_7/exppostnorm [0]) );
  AND2X1 U7157 ( .IN1(n5454), .IN2(n5442), .Q(
        \add_2_root_sub_1_root_fmul_0_0_0_0_7/add_321/carry [1]) );
  XOR2X1 U7158 ( .IN1(n5442), .IN2(n5454), .Q(
        \add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/A[0] ) );
  XNOR2X1 U7159 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/A[5] ), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/carry [5]), .Q(
        \fmul_0_0_0_0_6/exppostnorm [5]) );
  OR2X1 U7160 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/carry [4]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/A[4] ), .Q(
        \add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/carry [5]) );
  XNOR2X1 U7161 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/A[4] ), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/carry [4]), .Q(
        \fmul_0_0_0_0_6/exppostnorm [4]) );
  AND2X1 U7162 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/carry [3]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/A[3] ), .Q(
        \add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/carry [4]) );
  XOR2X1 U7163 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/carry [3]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/A[3] ), .Q(
        \fmul_0_0_0_0_6/exppostnorm [3]) );
  AND2X1 U7164 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/carry [2]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/A[2] ), .Q(
        \add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/carry [3]) );
  XOR2X1 U7165 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/carry [2]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/A[2] ), .Q(
        \fmul_0_0_0_0_6/exppostnorm [2]) );
  AND2X1 U7166 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/B[0] ), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/A[0] ), .Q(
        \add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/carry [1]) );
  XOR2X1 U7167 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/B[0] ), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/A[0] ), .Q(
        \fmul_0_0_0_0_6/exppostnorm [0]) );
  AND2X1 U7168 ( .IN1(n5526), .IN2(n5514), .Q(
        \add_2_root_sub_1_root_fmul_0_0_0_0_6/add_321/carry [1]) );
  XOR2X1 U7169 ( .IN1(n5514), .IN2(n5526), .Q(
        \add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/A[0] ) );
  XNOR2X1 U7170 ( .IN1(\fadd_0_0_0_0_5/newx_d1 [8]), .IN2(
        \fadd_0_0_0_0_5/sub_784/carry [4]), .Q(
        \fadd_0_0_0_0_5/exponentresultclose [4]) );
  OR2X1 U7171 ( .IN1(\fadd_0_0_0_0_5/sub_784/carry [3]), .IN2(
        \fadd_0_0_0_0_5/newx_d1 [7]), .Q(\fadd_0_0_0_0_5/sub_784/carry [4]) );
  XNOR2X1 U7172 ( .IN1(\fadd_0_0_0_0_5/newx_d1 [7]), .IN2(
        \fadd_0_0_0_0_5/sub_784/carry [3]), .Q(
        \fadd_0_0_0_0_5/exponentresultclose [3]) );
  OR2X1 U7173 ( .IN1(n14596), .IN2(\fadd_0_0_0_0_5/newx_d1 [4]), .Q(
        \fadd_0_0_0_0_5/sub_784/carry [1]) );
  XNOR2X1 U7174 ( .IN1(\fadd_0_0_0_0_5/newx_d1 [4]), .IN2(n14596), .Q(
        \fadd_0_0_0_0_5/exponentresultclose [0]) );
  XOR2X1 U7175 ( .IN1(
        \add_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [10]), .IN2(\fadd_0_0_0_0_5/resultbeforeround [10]), .Q(
        \fadd_0_0_0_0_5/resultrounded [10]) );
  XOR2X1 U7176 ( .IN1(n14229), .IN2(\fadd_0_0_0_0_5/add_859/carry [6]), .Q(
        \fadd_0_0_0_0_5/exponentresultfar1 [6]) );
  AND2X1 U7177 ( .IN1(
        \add_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [9]), .IN2(\fadd_0_0_0_0_5/resultbeforeround [9]), .Q(
        \add_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [10]) );
  XOR2X1 U7178 ( .IN1(
        \add_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [9]), .IN2(\fadd_0_0_0_0_5/resultbeforeround [9]), .Q(
        \fadd_0_0_0_0_5/resultrounded [9]) );
  AND2X1 U7179 ( .IN1(
        \add_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [8]), .IN2(\fadd_0_0_0_0_5/resultbeforeround [8]), .Q(
        \add_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [9]) );
  XOR2X1 U7180 ( .IN1(
        \add_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [8]), .IN2(\fadd_0_0_0_0_5/resultbeforeround [8]), .Q(
        \fadd_0_0_0_0_5/resultrounded [8]) );
  AND2X1 U7181 ( .IN1(
        \add_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [7]), .IN2(\fadd_0_0_0_0_5/resultbeforeround [7]), .Q(
        \add_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [8]) );
  XOR2X1 U7182 ( .IN1(
        \add_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [7]), .IN2(\fadd_0_0_0_0_5/resultbeforeround [7]), .Q(
        \fadd_0_0_0_0_5/resultrounded [7]) );
  AND2X1 U7183 ( .IN1(
        \add_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [6]), .IN2(\fadd_0_0_0_0_5/resultbeforeround [6]), .Q(
        \add_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [7]) );
  XOR2X1 U7184 ( .IN1(
        \add_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [6]), .IN2(\fadd_0_0_0_0_5/resultbeforeround [6]), .Q(
        \fadd_0_0_0_0_5/resultrounded [6]) );
  AND2X1 U7185 ( .IN1(
        \add_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [5]), .IN2(\fadd_0_0_0_0_5/resultbeforeround [5]), .Q(
        \add_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [6]) );
  XOR2X1 U7186 ( .IN1(
        \add_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [5]), .IN2(\fadd_0_0_0_0_5/resultbeforeround [5]), .Q(
        \fadd_0_0_0_0_5/resultrounded [5]) );
  AND2X1 U7187 ( .IN1(
        \add_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [4]), .IN2(\fadd_0_0_0_0_5/resultbeforeround [4]), .Q(
        \add_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [5]) );
  XOR2X1 U7188 ( .IN1(
        \add_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [4]), .IN2(\fadd_0_0_0_0_5/resultbeforeround [4]), .Q(
        \fadd_0_0_0_0_5/resultrounded [4]) );
  AND2X1 U7189 ( .IN1(
        \add_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [3]), .IN2(\fadd_0_0_0_0_5/resultbeforeround [3]), .Q(
        \add_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [4]) );
  XOR2X1 U7190 ( .IN1(
        \add_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [3]), .IN2(\fadd_0_0_0_0_5/resultbeforeround [3]), .Q(
        \fadd_0_0_0_0_5/resultrounded [3]) );
  AND2X1 U7191 ( .IN1(
        \add_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [2]), .IN2(\fadd_0_0_0_0_5/resultbeforeround [2]), .Q(
        \add_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [3]) );
  XOR2X1 U7192 ( .IN1(
        \add_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [2]), .IN2(\fadd_0_0_0_0_5/resultbeforeround [2]), .Q(
        \fadd_0_0_0_0_5/resultrounded [2]) );
  AND2X1 U7193 ( .IN1(
        \add_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [1]), .IN2(\fadd_0_0_0_0_5/resultbeforeround [1]), .Q(
        \add_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [2]) );
  XOR2X1 U7194 ( .IN1(
        \add_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [1]), .IN2(\fadd_0_0_0_0_5/resultbeforeround [1]), .Q(
        \fadd_0_0_0_0_5/resultrounded [1]) );
  AND2X1 U7195 ( .IN1(n14229), .IN2(\fadd_0_0_0_0_5/add_859/carry [5]), .Q(
        \fadd_0_0_0_0_5/add_859/carry [6]) );
  XOR2X1 U7196 ( .IN1(n14229), .IN2(\fadd_0_0_0_0_5/add_859/carry [5]), .Q(
        \fadd_0_0_0_0_5/exponentresultfar1 [5]) );
  AND2X1 U7197 ( .IN1(\fadd_0_0_0_0_5/expoperationsel[0] ), .IN2(
        \fadd_0_0_0_0_5/exponentresultfar0_d2 [0]), .Q(
        \fadd_0_0_0_0_5/add_859/carry [1]) );
  XOR2X1 U7198 ( .IN1(\fadd_0_0_0_0_5/expoperationsel[0] ), .IN2(
        \fadd_0_0_0_0_5/exponentresultfar0_d2 [0]), .Q(
        \fadd_0_0_0_0_5/exponentresultfar1 [0]) );
  AND2X1 U7199 ( .IN1(\fadd_0_0_0_0_5/round ), .IN2(
        \fadd_0_0_0_0_5/resultbeforeround [0]), .Q(
        \add_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [1]) );
  XOR2X1 U7200 ( .IN1(\fadd_0_0_0_0_5/round ), .IN2(
        \fadd_0_0_0_0_5/resultbeforeround [0]), .Q(
        \fadd_0_0_0_0_5/resultrounded [0]) );
  XOR2X1 U7201 ( .IN1(
        \add_1_root_fmul_0_0_0_0_5/roundingadder/add_57/carry [10]), .IN2(
        \fmul_0_0_0_0_5/roundingadder/x_1_d1 [10]), .Q(
        \fmul_0_0_0_0_5/expsigpostround [10]) );
  AND2X1 U7202 ( .IN1(
        \add_1_root_fmul_0_0_0_0_5/roundingadder/add_57/carry [9]), .IN2(
        \fmul_0_0_0_0_5/roundingadder/x_1_d1 [9]), .Q(
        \add_1_root_fmul_0_0_0_0_5/roundingadder/add_57/carry [10]) );
  XOR2X1 U7203 ( .IN1(
        \add_1_root_fmul_0_0_0_0_5/roundingadder/add_57/carry [9]), .IN2(
        \fmul_0_0_0_0_5/roundingadder/x_1_d1 [9]), .Q(
        \fmul_0_0_0_0_5/expsigpostround [9]) );
  AND2X1 U7204 ( .IN1(\fmul_0_0_0_0_5/roundingadder/x_1_d1 [8]), .IN2(
        \add_1_root_fmul_0_0_0_0_5/roundingadder/add_57/carry [8]), .Q(
        \add_1_root_fmul_0_0_0_0_5/roundingadder/add_57/carry [9]) );
  XOR2X1 U7205 ( .IN1(
        \add_1_root_fmul_0_0_0_0_5/roundingadder/add_57/carry [8]), .IN2(
        \fmul_0_0_0_0_5/roundingadder/x_1_d1 [8]), .Q(\U282/DATA2_8 ) );
  AND2X1 U7206 ( .IN1(\fmul_0_0_0_0_5/roundingadder/x_1_d1 [7]), .IN2(
        \add_1_root_fmul_0_0_0_0_5/roundingadder/add_57/carry [7]), .Q(
        \add_1_root_fmul_0_0_0_0_5/roundingadder/add_57/carry [8]) );
  XOR2X1 U7207 ( .IN1(
        \add_1_root_fmul_0_0_0_0_5/roundingadder/add_57/carry [7]), .IN2(
        \fmul_0_0_0_0_5/roundingadder/x_1_d1 [7]), .Q(\U282/DATA2_7 ) );
  AND2X1 U7208 ( .IN1(\fmul_0_0_0_0_5/roundingadder/x_1_d1 [6]), .IN2(
        \add_1_root_fmul_0_0_0_0_5/roundingadder/add_57/carry [6]), .Q(
        \add_1_root_fmul_0_0_0_0_5/roundingadder/add_57/carry [7]) );
  XOR2X1 U7209 ( .IN1(
        \add_1_root_fmul_0_0_0_0_5/roundingadder/add_57/carry [6]), .IN2(
        \fmul_0_0_0_0_5/roundingadder/x_1_d1 [6]), .Q(\U282/DATA2_6 ) );
  AND2X1 U7210 ( .IN1(\fmul_0_0_0_0_5/roundingadder/x_1_d1 [5]), .IN2(
        \add_1_root_fmul_0_0_0_0_5/roundingadder/add_57/carry [5]), .Q(
        \add_1_root_fmul_0_0_0_0_5/roundingadder/add_57/carry [6]) );
  XOR2X1 U7211 ( .IN1(
        \add_1_root_fmul_0_0_0_0_5/roundingadder/add_57/carry [5]), .IN2(
        \fmul_0_0_0_0_5/roundingadder/x_1_d1 [5]), .Q(\U282/DATA2_5 ) );
  AND2X1 U7212 ( .IN1(\fmul_0_0_0_0_5/roundingadder/x_1_d1 [4]), .IN2(
        \add_1_root_fmul_0_0_0_0_5/roundingadder/add_57/carry [4]), .Q(
        \add_1_root_fmul_0_0_0_0_5/roundingadder/add_57/carry [5]) );
  XOR2X1 U7213 ( .IN1(
        \add_1_root_fmul_0_0_0_0_5/roundingadder/add_57/carry [4]), .IN2(
        \fmul_0_0_0_0_5/roundingadder/x_1_d1 [4]), .Q(\U282/DATA2_4 ) );
  AND2X1 U7214 ( .IN1(\fmul_0_0_0_0_5/roundingadder/x_1_d1 [3]), .IN2(
        \add_1_root_fmul_0_0_0_0_5/roundingadder/add_57/carry [3]), .Q(
        \add_1_root_fmul_0_0_0_0_5/roundingadder/add_57/carry [4]) );
  XOR2X1 U7215 ( .IN1(
        \add_1_root_fmul_0_0_0_0_5/roundingadder/add_57/carry [3]), .IN2(
        \fmul_0_0_0_0_5/roundingadder/x_1_d1 [3]), .Q(\U282/DATA2_3 ) );
  AND2X1 U7216 ( .IN1(\fmul_0_0_0_0_5/roundingadder/x_1_d1 [2]), .IN2(
        \add_1_root_fmul_0_0_0_0_5/roundingadder/add_57/carry [2]), .Q(
        \add_1_root_fmul_0_0_0_0_5/roundingadder/add_57/carry [3]) );
  XOR2X1 U7217 ( .IN1(
        \add_1_root_fmul_0_0_0_0_5/roundingadder/add_57/carry [2]), .IN2(
        \fmul_0_0_0_0_5/roundingadder/x_1_d1 [2]), .Q(\U282/DATA2_2 ) );
  AND2X1 U7218 ( .IN1(\fmul_0_0_0_0_5/roundingadder/x_1_d1 [1]), .IN2(
        \add_1_root_fmul_0_0_0_0_5/roundingadder/add_57/carry [1]), .Q(
        \add_1_root_fmul_0_0_0_0_5/roundingadder/add_57/carry [2]) );
  XOR2X1 U7219 ( .IN1(
        \add_1_root_fmul_0_0_0_0_5/roundingadder/add_57/carry [1]), .IN2(
        \fmul_0_0_0_0_5/roundingadder/x_1_d1 [1]), .Q(\U282/DATA2_1 ) );
  AND2X1 U7220 ( .IN1(\fmul_0_0_0_0_5/roundingadder/n151_o[0] ), .IN2(
        \fmul_0_0_0_0_5/roundingadder/x_1_d1 [0]), .Q(
        \add_1_root_fmul_0_0_0_0_5/roundingadder/add_57/carry [1]) );
  XOR2X1 U7221 ( .IN1(\fmul_0_0_0_0_5/roundingadder/n151_o[0] ), .IN2(
        \fmul_0_0_0_0_5/roundingadder/x_1_d1 [0]), .Q(n13465) );
  XNOR2X1 U7222 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/A[5] ), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/carry [5]), .Q(
        \fmul_0_0_0_0_5/exppostnorm [5]) );
  OR2X1 U7223 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/carry [4]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/A[4] ), .Q(
        \add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/carry [5]) );
  XNOR2X1 U7224 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/A[4] ), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/carry [4]), .Q(
        \fmul_0_0_0_0_5/exppostnorm [4]) );
  AND2X1 U7225 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/carry [3]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/A[3] ), .Q(
        \add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/carry [4]) );
  XOR2X1 U7226 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/carry [3]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/A[3] ), .Q(
        \fmul_0_0_0_0_5/exppostnorm [3]) );
  AND2X1 U7227 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/carry [2]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/A[2] ), .Q(
        \add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/carry [3]) );
  XOR2X1 U7228 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/carry [2]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/A[2] ), .Q(
        \fmul_0_0_0_0_5/exppostnorm [2]) );
  AND2X1 U7229 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/B[0] ), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/A[0] ), .Q(
        \add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/carry [1]) );
  XOR2X1 U7230 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/B[0] ), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/A[0] ), .Q(
        \fmul_0_0_0_0_5/exppostnorm [0]) );
  AND2X1 U7231 ( .IN1(n5598), .IN2(n5586), .Q(
        \add_2_root_sub_1_root_fmul_0_0_0_0_5/add_321/carry [1]) );
  XOR2X1 U7232 ( .IN1(n5586), .IN2(n5598), .Q(
        \add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/A[0] ) );
  XNOR2X1 U7233 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/A[5] ), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/carry [5]), .Q(
        \fmul_0_0_0_0_4/exppostnorm [5]) );
  OR2X1 U7234 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/carry [4]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/A[4] ), .Q(
        \add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/carry [5]) );
  XNOR2X1 U7235 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/A[4] ), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/carry [4]), .Q(
        \fmul_0_0_0_0_4/exppostnorm [4]) );
  AND2X1 U7236 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/carry [3]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/A[3] ), .Q(
        \add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/carry [4]) );
  XOR2X1 U7237 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/carry [3]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/A[3] ), .Q(
        \fmul_0_0_0_0_4/exppostnorm [3]) );
  AND2X1 U7238 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/carry [2]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/A[2] ), .Q(
        \add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/carry [3]) );
  XOR2X1 U7239 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/carry [2]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/A[2] ), .Q(
        \fmul_0_0_0_0_4/exppostnorm [2]) );
  AND2X1 U7240 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/B[0] ), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/A[0] ), .Q(
        \add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/carry [1]) );
  XOR2X1 U7241 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/B[0] ), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/A[0] ), .Q(
        \fmul_0_0_0_0_4/exppostnorm [0]) );
  AND2X1 U7242 ( .IN1(n5670), .IN2(n5658), .Q(
        \add_2_root_sub_1_root_fmul_0_0_0_0_4/add_321/carry [1]) );
  XOR2X1 U7243 ( .IN1(n5658), .IN2(n5670), .Q(
        \add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/A[0] ) );
  XNOR2X1 U7244 ( .IN1(\fadd_0_0_0_0_2/newx_d1 [8]), .IN2(
        \fadd_0_0_0_0_2/sub_784/carry [4]), .Q(
        \fadd_0_0_0_0_2/exponentresultclose [4]) );
  OR2X1 U7245 ( .IN1(\fadd_0_0_0_0_2/sub_784/carry [3]), .IN2(
        \fadd_0_0_0_0_2/newx_d1 [7]), .Q(\fadd_0_0_0_0_2/sub_784/carry [4]) );
  XNOR2X1 U7246 ( .IN1(\fadd_0_0_0_0_2/newx_d1 [7]), .IN2(
        \fadd_0_0_0_0_2/sub_784/carry [3]), .Q(
        \fadd_0_0_0_0_2/exponentresultclose [3]) );
  OR2X1 U7247 ( .IN1(n14563), .IN2(\fadd_0_0_0_0_2/newx_d1 [4]), .Q(
        \fadd_0_0_0_0_2/sub_784/carry [1]) );
  XNOR2X1 U7248 ( .IN1(\fadd_0_0_0_0_2/newx_d1 [4]), .IN2(n14563), .Q(
        \fadd_0_0_0_0_2/exponentresultclose [0]) );
  XOR2X1 U7249 ( .IN1(
        \add_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [10]), .IN2(\fadd_0_0_0_0_2/resultbeforeround [10]), .Q(
        \fadd_0_0_0_0_2/resultrounded [10]) );
  XOR2X1 U7250 ( .IN1(n14226), .IN2(\fadd_0_0_0_0_2/add_859/carry [6]), .Q(
        \fadd_0_0_0_0_2/exponentresultfar1 [6]) );
  AND2X1 U7251 ( .IN1(
        \add_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [9]), .IN2(\fadd_0_0_0_0_2/resultbeforeround [9]), .Q(
        \add_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [10]) );
  AND2X1 U7252 ( .IN1(n14226), .IN2(\fadd_0_0_0_0_2/add_859/carry [5]), .Q(
        \fadd_0_0_0_0_2/add_859/carry [6]) );
  XOR2X1 U7253 ( .IN1(n14226), .IN2(\fadd_0_0_0_0_2/add_859/carry [5]), .Q(
        \fadd_0_0_0_0_2/exponentresultfar1 [5]) );
  AND2X1 U7254 ( .IN1(
        \add_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [8]), .IN2(\fadd_0_0_0_0_2/resultbeforeround [8]), .Q(
        \add_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [9]) );
  XOR2X1 U7255 ( .IN1(
        \add_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [8]), .IN2(\fadd_0_0_0_0_2/resultbeforeround [8]), .Q(
        \fadd_0_0_0_0_2/resultrounded [8]) );
  AND2X1 U7256 ( .IN1(
        \add_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [7]), .IN2(\fadd_0_0_0_0_2/resultbeforeround [7]), .Q(
        \add_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [8]) );
  XOR2X1 U7257 ( .IN1(
        \add_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [7]), .IN2(\fadd_0_0_0_0_2/resultbeforeround [7]), .Q(
        \fadd_0_0_0_0_2/resultrounded [7]) );
  AND2X1 U7258 ( .IN1(
        \add_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [6]), .IN2(\fadd_0_0_0_0_2/resultbeforeround [6]), .Q(
        \add_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [7]) );
  XOR2X1 U7259 ( .IN1(
        \add_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [6]), .IN2(\fadd_0_0_0_0_2/resultbeforeround [6]), .Q(
        \fadd_0_0_0_0_2/resultrounded [6]) );
  AND2X1 U7260 ( .IN1(
        \add_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [5]), .IN2(\fadd_0_0_0_0_2/resultbeforeround [5]), .Q(
        \add_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [6]) );
  XOR2X1 U7261 ( .IN1(
        \add_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [5]), .IN2(\fadd_0_0_0_0_2/resultbeforeround [5]), .Q(
        \fadd_0_0_0_0_2/resultrounded [5]) );
  AND2X1 U7262 ( .IN1(
        \add_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [4]), .IN2(\fadd_0_0_0_0_2/resultbeforeround [4]), .Q(
        \add_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [5]) );
  XOR2X1 U7263 ( .IN1(
        \add_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [4]), .IN2(\fadd_0_0_0_0_2/resultbeforeround [4]), .Q(
        \fadd_0_0_0_0_2/resultrounded [4]) );
  AND2X1 U7264 ( .IN1(
        \add_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [3]), .IN2(\fadd_0_0_0_0_2/resultbeforeround [3]), .Q(
        \add_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [4]) );
  XOR2X1 U7265 ( .IN1(
        \add_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [3]), .IN2(\fadd_0_0_0_0_2/resultbeforeround [3]), .Q(
        \fadd_0_0_0_0_2/resultrounded [3]) );
  AND2X1 U7266 ( .IN1(
        \add_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [2]), .IN2(\fadd_0_0_0_0_2/resultbeforeround [2]), .Q(
        \add_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [3]) );
  XOR2X1 U7267 ( .IN1(
        \add_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [2]), .IN2(\fadd_0_0_0_0_2/resultbeforeround [2]), .Q(
        \fadd_0_0_0_0_2/resultrounded [2]) );
  AND2X1 U7268 ( .IN1(
        \add_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [1]), .IN2(\fadd_0_0_0_0_2/resultbeforeround [1]), .Q(
        \add_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [2]) );
  XOR2X1 U7269 ( .IN1(
        \add_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [1]), .IN2(\fadd_0_0_0_0_2/resultbeforeround [1]), .Q(
        \fadd_0_0_0_0_2/resultrounded [1]) );
  AND2X1 U7270 ( .IN1(\fadd_0_0_0_0_2/round ), .IN2(
        \fadd_0_0_0_0_2/resultbeforeround [0]), .Q(
        \add_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [1]) );
  XOR2X1 U7271 ( .IN1(\fadd_0_0_0_0_2/round ), .IN2(
        \fadd_0_0_0_0_2/resultbeforeround [0]), .Q(
        \fadd_0_0_0_0_2/resultrounded [0]) );
  AND2X1 U7272 ( .IN1(\fadd_0_0_0_0_2/expoperationsel[0] ), .IN2(
        \fadd_0_0_0_0_2/exponentresultfar0_d2 [0]), .Q(
        \fadd_0_0_0_0_2/add_859/carry [1]) );
  XOR2X1 U7273 ( .IN1(\fadd_0_0_0_0_2/expoperationsel[0] ), .IN2(
        \fadd_0_0_0_0_2/exponentresultfar0_d2 [0]), .Q(
        \fadd_0_0_0_0_2/exponentresultfar1 [0]) );
  XNOR2X1 U7274 ( .IN1(\fadd_0_0_0_0_3/newx_d1 [8]), .IN2(
        \fadd_0_0_0_0_3/sub_784/carry [4]), .Q(
        \fadd_0_0_0_0_3/exponentresultclose [4]) );
  OR2X1 U7275 ( .IN1(\fadd_0_0_0_0_3/sub_784/carry [3]), .IN2(
        \fadd_0_0_0_0_3/newx_d1 [7]), .Q(\fadd_0_0_0_0_3/sub_784/carry [4]) );
  XNOR2X1 U7276 ( .IN1(\fadd_0_0_0_0_3/newx_d1 [7]), .IN2(
        \fadd_0_0_0_0_3/sub_784/carry [3]), .Q(
        \fadd_0_0_0_0_3/exponentresultclose [3]) );
  OR2X1 U7277 ( .IN1(n14574), .IN2(\fadd_0_0_0_0_3/newx_d1 [4]), .Q(
        \fadd_0_0_0_0_3/sub_784/carry [1]) );
  XNOR2X1 U7278 ( .IN1(\fadd_0_0_0_0_3/newx_d1 [4]), .IN2(n14574), .Q(
        \fadd_0_0_0_0_3/exponentresultclose [0]) );
  XOR2X1 U7279 ( .IN1(
        \add_1_root_fmul_0_0_0_0_2/roundingadder/add_57/carry [10]), .IN2(
        \fmul_0_0_0_0_2/roundingadder/x_1_d1 [10]), .Q(
        \fmul_0_0_0_0_2/expsigpostround [10]) );
  AND2X1 U7280 ( .IN1(
        \add_1_root_fmul_0_0_0_0_2/roundingadder/add_57/carry [9]), .IN2(
        \fmul_0_0_0_0_2/roundingadder/x_1_d1 [9]), .Q(
        \add_1_root_fmul_0_0_0_0_2/roundingadder/add_57/carry [10]) );
  XOR2X1 U7281 ( .IN1(
        \add_1_root_fmul_0_0_0_0_2/roundingadder/add_57/carry [9]), .IN2(
        \fmul_0_0_0_0_2/roundingadder/x_1_d1 [9]), .Q(
        \fmul_0_0_0_0_2/expsigpostround [9]) );
  AND2X1 U7282 ( .IN1(\fmul_0_0_0_0_2/roundingadder/x_1_d1 [8]), .IN2(
        \add_1_root_fmul_0_0_0_0_2/roundingadder/add_57/carry [8]), .Q(
        \add_1_root_fmul_0_0_0_0_2/roundingadder/add_57/carry [9]) );
  XOR2X1 U7283 ( .IN1(
        \add_1_root_fmul_0_0_0_0_2/roundingadder/add_57/carry [8]), .IN2(
        \fmul_0_0_0_0_2/roundingadder/x_1_d1 [8]), .Q(\U450/DATA2_8 ) );
  AND2X1 U7284 ( .IN1(\fmul_0_0_0_0_2/roundingadder/x_1_d1 [7]), .IN2(
        \add_1_root_fmul_0_0_0_0_2/roundingadder/add_57/carry [7]), .Q(
        \add_1_root_fmul_0_0_0_0_2/roundingadder/add_57/carry [8]) );
  XOR2X1 U7285 ( .IN1(
        \add_1_root_fmul_0_0_0_0_2/roundingadder/add_57/carry [7]), .IN2(
        \fmul_0_0_0_0_2/roundingadder/x_1_d1 [7]), .Q(\U450/DATA2_7 ) );
  AND2X1 U7286 ( .IN1(\fmul_0_0_0_0_2/roundingadder/x_1_d1 [6]), .IN2(
        \add_1_root_fmul_0_0_0_0_2/roundingadder/add_57/carry [6]), .Q(
        \add_1_root_fmul_0_0_0_0_2/roundingadder/add_57/carry [7]) );
  XOR2X1 U7287 ( .IN1(
        \add_1_root_fmul_0_0_0_0_2/roundingadder/add_57/carry [6]), .IN2(
        \fmul_0_0_0_0_2/roundingadder/x_1_d1 [6]), .Q(\U450/DATA2_6 ) );
  AND2X1 U7288 ( .IN1(\fmul_0_0_0_0_2/roundingadder/x_1_d1 [5]), .IN2(
        \add_1_root_fmul_0_0_0_0_2/roundingadder/add_57/carry [5]), .Q(
        \add_1_root_fmul_0_0_0_0_2/roundingadder/add_57/carry [6]) );
  XOR2X1 U7289 ( .IN1(
        \add_1_root_fmul_0_0_0_0_2/roundingadder/add_57/carry [5]), .IN2(
        \fmul_0_0_0_0_2/roundingadder/x_1_d1 [5]), .Q(\U450/DATA2_5 ) );
  AND2X1 U7290 ( .IN1(\fmul_0_0_0_0_2/roundingadder/x_1_d1 [4]), .IN2(
        \add_1_root_fmul_0_0_0_0_2/roundingadder/add_57/carry [4]), .Q(
        \add_1_root_fmul_0_0_0_0_2/roundingadder/add_57/carry [5]) );
  XOR2X1 U7291 ( .IN1(
        \add_1_root_fmul_0_0_0_0_2/roundingadder/add_57/carry [4]), .IN2(
        \fmul_0_0_0_0_2/roundingadder/x_1_d1 [4]), .Q(\U450/DATA2_4 ) );
  AND2X1 U7292 ( .IN1(\fmul_0_0_0_0_2/roundingadder/x_1_d1 [3]), .IN2(
        \add_1_root_fmul_0_0_0_0_2/roundingadder/add_57/carry [3]), .Q(
        \add_1_root_fmul_0_0_0_0_2/roundingadder/add_57/carry [4]) );
  XOR2X1 U7293 ( .IN1(
        \add_1_root_fmul_0_0_0_0_2/roundingadder/add_57/carry [3]), .IN2(
        \fmul_0_0_0_0_2/roundingadder/x_1_d1 [3]), .Q(\U450/DATA2_3 ) );
  AND2X1 U7294 ( .IN1(\fmul_0_0_0_0_2/roundingadder/x_1_d1 [2]), .IN2(
        \add_1_root_fmul_0_0_0_0_2/roundingadder/add_57/carry [2]), .Q(
        \add_1_root_fmul_0_0_0_0_2/roundingadder/add_57/carry [3]) );
  XOR2X1 U7295 ( .IN1(
        \add_1_root_fmul_0_0_0_0_2/roundingadder/add_57/carry [2]), .IN2(
        \fmul_0_0_0_0_2/roundingadder/x_1_d1 [2]), .Q(\U450/DATA2_2 ) );
  AND2X1 U7296 ( .IN1(\fmul_0_0_0_0_2/roundingadder/x_1_d1 [1]), .IN2(
        \add_1_root_fmul_0_0_0_0_2/roundingadder/add_57/carry [1]), .Q(
        \add_1_root_fmul_0_0_0_0_2/roundingadder/add_57/carry [2]) );
  XOR2X1 U7297 ( .IN1(
        \add_1_root_fmul_0_0_0_0_2/roundingadder/add_57/carry [1]), .IN2(
        \fmul_0_0_0_0_2/roundingadder/x_1_d1 [1]), .Q(\U450/DATA2_1 ) );
  AND2X1 U7298 ( .IN1(\fmul_0_0_0_0_2/roundingadder/x_1_d1 [0]), .IN2(
        \fmul_0_0_0_0_2/roundingadder/n151_o[0] ), .Q(
        \add_1_root_fmul_0_0_0_0_2/roundingadder/add_57/carry [1]) );
  XOR2X1 U7299 ( .IN1(\fmul_0_0_0_0_2/roundingadder/n151_o[0] ), .IN2(
        \fmul_0_0_0_0_2/roundingadder/x_1_d1 [0]), .Q(\U450/DATA2_0 ) );
  XOR2X1 U7300 ( .IN1(
        \add_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [10]), .IN2(\fadd_0_0_0_0_3/resultbeforeround [10]), .Q(
        \fadd_0_0_0_0_3/resultrounded [10]) );
  XOR2X1 U7301 ( .IN1(n14227), .IN2(\fadd_0_0_0_0_3/add_859/carry [6]), .Q(
        \fadd_0_0_0_0_3/exponentresultfar1 [6]) );
  AND2X1 U7302 ( .IN1(
        \add_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [9]), .IN2(\fadd_0_0_0_0_3/resultbeforeround [9]), .Q(
        \add_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [10]) );
  XOR2X1 U7303 ( .IN1(
        \add_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [9]), .IN2(\fadd_0_0_0_0_3/resultbeforeround [9]), .Q(
        \fadd_0_0_0_0_3/resultrounded [9]) );
  AND2X1 U7304 ( .IN1(
        \add_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [8]), .IN2(\fadd_0_0_0_0_3/resultbeforeround [8]), .Q(
        \add_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [9]) );
  XOR2X1 U7305 ( .IN1(
        \add_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [8]), .IN2(\fadd_0_0_0_0_3/resultbeforeround [8]), .Q(
        \fadd_0_0_0_0_3/resultrounded [8]) );
  AND2X1 U7306 ( .IN1(
        \add_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [7]), .IN2(\fadd_0_0_0_0_3/resultbeforeround [7]), .Q(
        \add_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [8]) );
  XOR2X1 U7307 ( .IN1(
        \add_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [7]), .IN2(\fadd_0_0_0_0_3/resultbeforeround [7]), .Q(
        \fadd_0_0_0_0_3/resultrounded [7]) );
  AND2X1 U7308 ( .IN1(
        \add_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [6]), .IN2(\fadd_0_0_0_0_3/resultbeforeround [6]), .Q(
        \add_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [7]) );
  XOR2X1 U7309 ( .IN1(
        \add_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [6]), .IN2(\fadd_0_0_0_0_3/resultbeforeround [6]), .Q(
        \fadd_0_0_0_0_3/resultrounded [6]) );
  AND2X1 U7310 ( .IN1(
        \add_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [5]), .IN2(\fadd_0_0_0_0_3/resultbeforeround [5]), .Q(
        \add_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [6]) );
  XOR2X1 U7311 ( .IN1(
        \add_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [5]), .IN2(\fadd_0_0_0_0_3/resultbeforeround [5]), .Q(
        \fadd_0_0_0_0_3/resultrounded [5]) );
  AND2X1 U7312 ( .IN1(
        \add_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [4]), .IN2(\fadd_0_0_0_0_3/resultbeforeround [4]), .Q(
        \add_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [5]) );
  XOR2X1 U7313 ( .IN1(
        \add_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [4]), .IN2(\fadd_0_0_0_0_3/resultbeforeround [4]), .Q(
        \fadd_0_0_0_0_3/resultrounded [4]) );
  AND2X1 U7314 ( .IN1(
        \add_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [3]), .IN2(\fadd_0_0_0_0_3/resultbeforeround [3]), .Q(
        \add_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [4]) );
  XOR2X1 U7315 ( .IN1(
        \add_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [3]), .IN2(\fadd_0_0_0_0_3/resultbeforeround [3]), .Q(
        \fadd_0_0_0_0_3/resultrounded [3]) );
  AND2X1 U7316 ( .IN1(
        \add_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [2]), .IN2(\fadd_0_0_0_0_3/resultbeforeround [2]), .Q(
        \add_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [3]) );
  XOR2X1 U7317 ( .IN1(
        \add_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [2]), .IN2(\fadd_0_0_0_0_3/resultbeforeround [2]), .Q(
        \fadd_0_0_0_0_3/resultrounded [2]) );
  AND2X1 U7318 ( .IN1(
        \add_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [1]), .IN2(\fadd_0_0_0_0_3/resultbeforeround [1]), .Q(
        \add_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [2]) );
  XOR2X1 U7319 ( .IN1(
        \add_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [1]), .IN2(\fadd_0_0_0_0_3/resultbeforeround [1]), .Q(
        \fadd_0_0_0_0_3/resultrounded [1]) );
  AND2X1 U7320 ( .IN1(\fadd_0_0_0_0_3/round ), .IN2(
        \fadd_0_0_0_0_3/resultbeforeround [0]), .Q(
        \add_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [1]) );
  XOR2X1 U7321 ( .IN1(\fadd_0_0_0_0_3/round ), .IN2(
        \fadd_0_0_0_0_3/resultbeforeround [0]), .Q(
        \fadd_0_0_0_0_3/resultrounded [0]) );
  AND2X1 U7322 ( .IN1(n14227), .IN2(\fadd_0_0_0_0_3/add_859/carry [5]), .Q(
        \fadd_0_0_0_0_3/add_859/carry [6]) );
  XOR2X1 U7323 ( .IN1(n14227), .IN2(\fadd_0_0_0_0_3/add_859/carry [5]), .Q(
        \fadd_0_0_0_0_3/exponentresultfar1 [5]) );
  AND2X1 U7324 ( .IN1(\fadd_0_0_0_0_3/expoperationsel[0] ), .IN2(
        \fadd_0_0_0_0_3/exponentresultfar0_d2 [0]), .Q(
        \fadd_0_0_0_0_3/add_859/carry [1]) );
  XOR2X1 U7325 ( .IN1(\fadd_0_0_0_0_3/expoperationsel[0] ), .IN2(
        \fadd_0_0_0_0_3/exponentresultfar0_d2 [0]), .Q(
        \fadd_0_0_0_0_3/exponentresultfar1 [0]) );
  XOR2X1 U7326 ( .IN1(
        \add_1_root_fmul_0_0_0_0_3/roundingadder/add_57/carry [10]), .IN2(
        \fmul_0_0_0_0_3/roundingadder/x_1_d1 [10]), .Q(
        \fmul_0_0_0_0_3/expsigpostround [10]) );
  AND2X1 U7327 ( .IN1(
        \add_1_root_fmul_0_0_0_0_3/roundingadder/add_57/carry [9]), .IN2(
        \fmul_0_0_0_0_3/roundingadder/x_1_d1 [9]), .Q(
        \add_1_root_fmul_0_0_0_0_3/roundingadder/add_57/carry [10]) );
  XOR2X1 U7328 ( .IN1(
        \add_1_root_fmul_0_0_0_0_3/roundingadder/add_57/carry [9]), .IN2(
        \fmul_0_0_0_0_3/roundingadder/x_1_d1 [9]), .Q(
        \fmul_0_0_0_0_3/expsigpostround [9]) );
  AND2X1 U7329 ( .IN1(\fmul_0_0_0_0_3/roundingadder/x_1_d1 [8]), .IN2(
        \add_1_root_fmul_0_0_0_0_3/roundingadder/add_57/carry [8]), .Q(
        \add_1_root_fmul_0_0_0_0_3/roundingadder/add_57/carry [9]) );
  XOR2X1 U7330 ( .IN1(
        \add_1_root_fmul_0_0_0_0_3/roundingadder/add_57/carry [8]), .IN2(
        \fmul_0_0_0_0_3/roundingadder/x_1_d1 [8]), .Q(\U394/DATA2_8 ) );
  AND2X1 U7331 ( .IN1(\fmul_0_0_0_0_3/roundingadder/x_1_d1 [7]), .IN2(
        \add_1_root_fmul_0_0_0_0_3/roundingadder/add_57/carry [7]), .Q(
        \add_1_root_fmul_0_0_0_0_3/roundingadder/add_57/carry [8]) );
  XOR2X1 U7332 ( .IN1(
        \add_1_root_fmul_0_0_0_0_3/roundingadder/add_57/carry [7]), .IN2(
        \fmul_0_0_0_0_3/roundingadder/x_1_d1 [7]), .Q(\U394/DATA2_7 ) );
  AND2X1 U7333 ( .IN1(\fmul_0_0_0_0_3/roundingadder/x_1_d1 [6]), .IN2(
        \add_1_root_fmul_0_0_0_0_3/roundingadder/add_57/carry [6]), .Q(
        \add_1_root_fmul_0_0_0_0_3/roundingadder/add_57/carry [7]) );
  XOR2X1 U7334 ( .IN1(
        \add_1_root_fmul_0_0_0_0_3/roundingadder/add_57/carry [6]), .IN2(
        \fmul_0_0_0_0_3/roundingadder/x_1_d1 [6]), .Q(\U394/DATA2_6 ) );
  AND2X1 U7335 ( .IN1(\fmul_0_0_0_0_3/roundingadder/x_1_d1 [5]), .IN2(
        \add_1_root_fmul_0_0_0_0_3/roundingadder/add_57/carry [5]), .Q(
        \add_1_root_fmul_0_0_0_0_3/roundingadder/add_57/carry [6]) );
  XOR2X1 U7336 ( .IN1(
        \add_1_root_fmul_0_0_0_0_3/roundingadder/add_57/carry [5]), .IN2(
        \fmul_0_0_0_0_3/roundingadder/x_1_d1 [5]), .Q(\U394/DATA2_5 ) );
  AND2X1 U7337 ( .IN1(\fmul_0_0_0_0_3/roundingadder/x_1_d1 [4]), .IN2(
        \add_1_root_fmul_0_0_0_0_3/roundingadder/add_57/carry [4]), .Q(
        \add_1_root_fmul_0_0_0_0_3/roundingadder/add_57/carry [5]) );
  XOR2X1 U7338 ( .IN1(
        \add_1_root_fmul_0_0_0_0_3/roundingadder/add_57/carry [4]), .IN2(
        \fmul_0_0_0_0_3/roundingadder/x_1_d1 [4]), .Q(\U394/DATA2_4 ) );
  AND2X1 U7339 ( .IN1(\fmul_0_0_0_0_3/roundingadder/x_1_d1 [3]), .IN2(
        \add_1_root_fmul_0_0_0_0_3/roundingadder/add_57/carry [3]), .Q(
        \add_1_root_fmul_0_0_0_0_3/roundingadder/add_57/carry [4]) );
  XOR2X1 U7340 ( .IN1(
        \add_1_root_fmul_0_0_0_0_3/roundingadder/add_57/carry [3]), .IN2(
        \fmul_0_0_0_0_3/roundingadder/x_1_d1 [3]), .Q(\U394/DATA2_3 ) );
  AND2X1 U7341 ( .IN1(\fmul_0_0_0_0_3/roundingadder/x_1_d1 [2]), .IN2(
        \add_1_root_fmul_0_0_0_0_3/roundingadder/add_57/carry [2]), .Q(
        \add_1_root_fmul_0_0_0_0_3/roundingadder/add_57/carry [3]) );
  XOR2X1 U7342 ( .IN1(
        \add_1_root_fmul_0_0_0_0_3/roundingadder/add_57/carry [2]), .IN2(
        \fmul_0_0_0_0_3/roundingadder/x_1_d1 [2]), .Q(\U394/DATA2_2 ) );
  AND2X1 U7343 ( .IN1(\fmul_0_0_0_0_3/roundingadder/x_1_d1 [1]), .IN2(
        \add_1_root_fmul_0_0_0_0_3/roundingadder/add_57/carry [1]), .Q(
        \add_1_root_fmul_0_0_0_0_3/roundingadder/add_57/carry [2]) );
  XOR2X1 U7344 ( .IN1(
        \add_1_root_fmul_0_0_0_0_3/roundingadder/add_57/carry [1]), .IN2(
        \fmul_0_0_0_0_3/roundingadder/x_1_d1 [1]), .Q(\U394/DATA2_1 ) );
  AND2X1 U7345 ( .IN1(\fmul_0_0_0_0_3/roundingadder/x_1_d1 [0]), .IN2(
        \fmul_0_0_0_0_3/roundingadder/n151_o[0] ), .Q(
        \add_1_root_fmul_0_0_0_0_3/roundingadder/add_57/carry [1]) );
  XOR2X1 U7346 ( .IN1(\fmul_0_0_0_0_3/roundingadder/n151_o[0] ), .IN2(
        \fmul_0_0_0_0_3/roundingadder/x_1_d1 [0]), .Q(\U394/DATA2_0 ) );
  XNOR2X1 U7347 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/A[5] ), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/carry [5]), .Q(
        \fmul_0_0_0_0_3/exppostnorm [5]) );
  OR2X1 U7348 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/carry [4]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/A[4] ), .Q(
        \add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/carry [5]) );
  XNOR2X1 U7349 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/A[4] ), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/carry [4]), .Q(
        \fmul_0_0_0_0_3/exppostnorm [4]) );
  AND2X1 U7350 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/carry [3]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/A[3] ), .Q(
        \add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/carry [4]) );
  XOR2X1 U7351 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/carry [3]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/A[3] ), .Q(
        \fmul_0_0_0_0_3/exppostnorm [3]) );
  AND2X1 U7352 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/carry [2]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/A[2] ), .Q(
        \add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/carry [3]) );
  XOR2X1 U7353 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/carry [2]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/A[2] ), .Q(
        \fmul_0_0_0_0_3/exppostnorm [2]) );
  AND2X1 U7354 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/B[0] ), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/A[0] ), .Q(
        \add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/carry [1]) );
  XOR2X1 U7355 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/B[0] ), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/A[0] ), .Q(
        \fmul_0_0_0_0_3/exppostnorm [0]) );
  AND2X1 U7356 ( .IN1(n5742), .IN2(n5730), .Q(
        \add_2_root_sub_1_root_fmul_0_0_0_0_3/add_321/carry [1]) );
  XOR2X1 U7357 ( .IN1(n5730), .IN2(n5742), .Q(
        \add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/A[0] ) );
  XNOR2X1 U7358 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/A[5] ), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/carry [5]), .Q(
        \fmul_0_0_0_0_2/exppostnorm [5]) );
  OR2X1 U7359 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/carry [4]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/A[4] ), .Q(
        \add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/carry [5]) );
  XNOR2X1 U7360 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/A[4] ), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/carry [4]), .Q(
        \fmul_0_0_0_0_2/exppostnorm [4]) );
  AND2X1 U7361 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/carry [3]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/A[3] ), .Q(
        \add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/carry [4]) );
  XOR2X1 U7362 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/carry [3]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/A[3] ), .Q(
        \fmul_0_0_0_0_2/exppostnorm [3]) );
  AND2X1 U7363 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/carry [2]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/A[2] ), .Q(
        \add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/carry [3]) );
  XOR2X1 U7364 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/carry [2]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/A[2] ), .Q(
        \fmul_0_0_0_0_2/exppostnorm [2]) );
  AND2X1 U7365 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/B[0] ), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/A[0] ), .Q(
        \add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/carry [1]) );
  XOR2X1 U7366 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/B[0] ), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/A[0] ), .Q(
        \fmul_0_0_0_0_2/exppostnorm [0]) );
  AND2X1 U7367 ( .IN1(n5814), .IN2(n5802), .Q(
        \add_2_root_sub_1_root_fmul_0_0_0_0_2/add_321/carry [1]) );
  XOR2X1 U7368 ( .IN1(n5802), .IN2(n5814), .Q(
        \add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/A[0] ) );
  XNOR2X1 U7369 ( .IN1(\fadd_0_0_0_0_1/newx_d1 [8]), .IN2(
        \fadd_0_0_0_0_1/sub_784/carry [4]), .Q(
        \fadd_0_0_0_0_1/exponentresultclose [4]) );
  OR2X1 U7370 ( .IN1(\fadd_0_0_0_0_1/sub_784/carry [3]), .IN2(
        \fadd_0_0_0_0_1/newx_d1 [7]), .Q(\fadd_0_0_0_0_1/sub_784/carry [4]) );
  XNOR2X1 U7371 ( .IN1(\fadd_0_0_0_0_1/newx_d1 [7]), .IN2(
        \fadd_0_0_0_0_1/sub_784/carry [3]), .Q(
        \fadd_0_0_0_0_1/exponentresultclose [3]) );
  OR2X1 U7372 ( .IN1(n14552), .IN2(\fadd_0_0_0_0_1/newx_d1 [4]), .Q(
        \fadd_0_0_0_0_1/sub_784/carry [1]) );
  XNOR2X1 U7373 ( .IN1(\fadd_0_0_0_0_1/newx_d1 [4]), .IN2(n14552), .Q(
        \fadd_0_0_0_0_1/exponentresultclose [0]) );
  XOR2X1 U7374 ( .IN1(
        \add_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [10]), .IN2(\fadd_0_0_0_0_1/resultbeforeround [10]), .Q(
        \fadd_0_0_0_0_1/resultrounded [10]) );
  XOR2X1 U7375 ( .IN1(\fadd_0_0_0_0_1/add_859/B[1] ), .IN2(
        \fadd_0_0_0_0_1/add_859/carry [6]), .Q(
        \fadd_0_0_0_0_1/exponentresultfar1 [6]) );
  AND2X1 U7376 ( .IN1(
        \add_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [9]), .IN2(\fadd_0_0_0_0_1/resultbeforeround [9]), .Q(
        \add_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [10]) );
  XOR2X1 U7377 ( .IN1(
        \add_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [9]), .IN2(\fadd_0_0_0_0_1/resultbeforeround [9]), .Q(
        \fadd_0_0_0_0_1/resultrounded [9]) );
  AND2X1 U7378 ( .IN1(
        \add_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [8]), .IN2(\fadd_0_0_0_0_1/resultbeforeround [8]), .Q(
        \add_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [9]) );
  XOR2X1 U7379 ( .IN1(
        \add_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [8]), .IN2(\fadd_0_0_0_0_1/resultbeforeround [8]), .Q(
        \fadd_0_0_0_0_1/resultrounded [8]) );
  AND2X1 U7380 ( .IN1(
        \add_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [7]), .IN2(\fadd_0_0_0_0_1/resultbeforeround [7]), .Q(
        \add_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [8]) );
  XOR2X1 U7381 ( .IN1(
        \add_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [7]), .IN2(\fadd_0_0_0_0_1/resultbeforeround [7]), .Q(
        \fadd_0_0_0_0_1/resultrounded [7]) );
  AND2X1 U7382 ( .IN1(
        \add_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [6]), .IN2(\fadd_0_0_0_0_1/resultbeforeround [6]), .Q(
        \add_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [7]) );
  XOR2X1 U7383 ( .IN1(
        \add_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [6]), .IN2(\fadd_0_0_0_0_1/resultbeforeround [6]), .Q(
        \fadd_0_0_0_0_1/resultrounded [6]) );
  AND2X1 U7384 ( .IN1(
        \add_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [5]), .IN2(\fadd_0_0_0_0_1/resultbeforeround [5]), .Q(
        \add_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [6]) );
  XOR2X1 U7385 ( .IN1(
        \add_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [5]), .IN2(\fadd_0_0_0_0_1/resultbeforeround [5]), .Q(
        \fadd_0_0_0_0_1/resultrounded [5]) );
  AND2X1 U7386 ( .IN1(
        \add_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [4]), .IN2(\fadd_0_0_0_0_1/resultbeforeround [4]), .Q(
        \add_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [5]) );
  XOR2X1 U7387 ( .IN1(
        \add_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [4]), .IN2(\fadd_0_0_0_0_1/resultbeforeround [4]), .Q(
        \fadd_0_0_0_0_1/resultrounded [4]) );
  AND2X1 U7388 ( .IN1(
        \add_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [3]), .IN2(\fadd_0_0_0_0_1/resultbeforeround [3]), .Q(
        \add_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [4]) );
  XOR2X1 U7389 ( .IN1(
        \add_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [3]), .IN2(\fadd_0_0_0_0_1/resultbeforeround [3]), .Q(
        \fadd_0_0_0_0_1/resultrounded [3]) );
  AND2X1 U7390 ( .IN1(
        \add_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [2]), .IN2(\fadd_0_0_0_0_1/resultbeforeround [2]), .Q(
        \add_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [3]) );
  XOR2X1 U7391 ( .IN1(
        \add_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [2]), .IN2(\fadd_0_0_0_0_1/resultbeforeround [2]), .Q(
        \fadd_0_0_0_0_1/resultrounded [2]) );
  AND2X1 U7392 ( .IN1(
        \add_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [1]), .IN2(\fadd_0_0_0_0_1/resultbeforeround [1]), .Q(
        \add_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [2]) );
  XOR2X1 U7393 ( .IN1(
        \add_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [1]), .IN2(\fadd_0_0_0_0_1/resultbeforeround [1]), .Q(
        \fadd_0_0_0_0_1/resultrounded [1]) );
  AND2X1 U7394 ( .IN1(\fadd_0_0_0_0_1/round ), .IN2(
        \fadd_0_0_0_0_1/resultbeforeround [0]), .Q(
        \add_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_finalroundadd/add_21/carry [1]) );
  XOR2X1 U7395 ( .IN1(\fadd_0_0_0_0_1/round ), .IN2(
        \fadd_0_0_0_0_1/resultbeforeround [0]), .Q(
        \fadd_0_0_0_0_1/resultrounded [0]) );
  AND2X1 U7396 ( .IN1(\fadd_0_0_0_0_1/add_859/B[1] ), .IN2(
        \fadd_0_0_0_0_1/add_859/carry [5]), .Q(
        \fadd_0_0_0_0_1/add_859/carry [6]) );
  XOR2X1 U7397 ( .IN1(\fadd_0_0_0_0_1/add_859/B[1] ), .IN2(
        \fadd_0_0_0_0_1/add_859/carry [5]), .Q(
        \fadd_0_0_0_0_1/exponentresultfar1 [5]) );
  AND2X1 U7398 ( .IN1(\fadd_0_0_0_0_1/expoperationsel[0] ), .IN2(
        \fadd_0_0_0_0_1/exponentresultfar0_d2 [0]), .Q(
        \fadd_0_0_0_0_1/add_859/carry [1]) );
  XOR2X1 U7399 ( .IN1(\fadd_0_0_0_0_1/expoperationsel[0] ), .IN2(
        \fadd_0_0_0_0_1/exponentresultfar0_d2 [0]), .Q(
        \fadd_0_0_0_0_1/exponentresultfar1 [0]) );
  XOR2X1 U7400 ( .IN1(
        \add_1_root_fmul_0_0_0_0_1/roundingadder/add_57/carry [10]), .IN2(
        \fmul_0_0_0_0_1/roundingadder/x_1_d1 [10]), .Q(
        \fmul_0_0_0_0_1/expsigpostround [10]) );
  AND2X1 U7401 ( .IN1(
        \add_1_root_fmul_0_0_0_0_1/roundingadder/add_57/carry [9]), .IN2(
        \fmul_0_0_0_0_1/roundingadder/x_1_d1 [9]), .Q(
        \add_1_root_fmul_0_0_0_0_1/roundingadder/add_57/carry [10]) );
  XOR2X1 U7402 ( .IN1(
        \add_1_root_fmul_0_0_0_0_1/roundingadder/add_57/carry [9]), .IN2(
        \fmul_0_0_0_0_1/roundingadder/x_1_d1 [9]), .Q(
        \fmul_0_0_0_0_1/expsigpostround [9]) );
  AND2X1 U7403 ( .IN1(\fmul_0_0_0_0_1/roundingadder/x_1_d1 [8]), .IN2(
        \add_1_root_fmul_0_0_0_0_1/roundingadder/add_57/carry [8]), .Q(
        \add_1_root_fmul_0_0_0_0_1/roundingadder/add_57/carry [9]) );
  XOR2X1 U7404 ( .IN1(
        \add_1_root_fmul_0_0_0_0_1/roundingadder/add_57/carry [8]), .IN2(
        \fmul_0_0_0_0_1/roundingadder/x_1_d1 [8]), .Q(\U503/DATA2_8 ) );
  AND2X1 U7405 ( .IN1(\fmul_0_0_0_0_1/roundingadder/x_1_d1 [7]), .IN2(
        \add_1_root_fmul_0_0_0_0_1/roundingadder/add_57/carry [7]), .Q(
        \add_1_root_fmul_0_0_0_0_1/roundingadder/add_57/carry [8]) );
  XOR2X1 U7406 ( .IN1(
        \add_1_root_fmul_0_0_0_0_1/roundingadder/add_57/carry [7]), .IN2(
        \fmul_0_0_0_0_1/roundingadder/x_1_d1 [7]), .Q(\U503/DATA2_7 ) );
  AND2X1 U7407 ( .IN1(\fmul_0_0_0_0_1/roundingadder/x_1_d1 [6]), .IN2(
        \add_1_root_fmul_0_0_0_0_1/roundingadder/add_57/carry [6]), .Q(
        \add_1_root_fmul_0_0_0_0_1/roundingadder/add_57/carry [7]) );
  XOR2X1 U7408 ( .IN1(
        \add_1_root_fmul_0_0_0_0_1/roundingadder/add_57/carry [6]), .IN2(
        \fmul_0_0_0_0_1/roundingadder/x_1_d1 [6]), .Q(\U503/DATA2_6 ) );
  AND2X1 U7409 ( .IN1(\fmul_0_0_0_0_1/roundingadder/x_1_d1 [5]), .IN2(
        \add_1_root_fmul_0_0_0_0_1/roundingadder/add_57/carry [5]), .Q(
        \add_1_root_fmul_0_0_0_0_1/roundingadder/add_57/carry [6]) );
  XOR2X1 U7410 ( .IN1(
        \add_1_root_fmul_0_0_0_0_1/roundingadder/add_57/carry [5]), .IN2(
        \fmul_0_0_0_0_1/roundingadder/x_1_d1 [5]), .Q(\U503/DATA2_5 ) );
  AND2X1 U7411 ( .IN1(\fmul_0_0_0_0_1/roundingadder/x_1_d1 [4]), .IN2(
        \add_1_root_fmul_0_0_0_0_1/roundingadder/add_57/carry [4]), .Q(
        \add_1_root_fmul_0_0_0_0_1/roundingadder/add_57/carry [5]) );
  XOR2X1 U7412 ( .IN1(
        \add_1_root_fmul_0_0_0_0_1/roundingadder/add_57/carry [4]), .IN2(
        \fmul_0_0_0_0_1/roundingadder/x_1_d1 [4]), .Q(\U503/DATA2_4 ) );
  AND2X1 U7413 ( .IN1(\fmul_0_0_0_0_1/roundingadder/x_1_d1 [3]), .IN2(
        \add_1_root_fmul_0_0_0_0_1/roundingadder/add_57/carry [3]), .Q(
        \add_1_root_fmul_0_0_0_0_1/roundingadder/add_57/carry [4]) );
  XOR2X1 U7414 ( .IN1(
        \add_1_root_fmul_0_0_0_0_1/roundingadder/add_57/carry [3]), .IN2(
        \fmul_0_0_0_0_1/roundingadder/x_1_d1 [3]), .Q(\U503/DATA2_3 ) );
  AND2X1 U7415 ( .IN1(\fmul_0_0_0_0_1/roundingadder/x_1_d1 [2]), .IN2(
        \add_1_root_fmul_0_0_0_0_1/roundingadder/add_57/carry [2]), .Q(
        \add_1_root_fmul_0_0_0_0_1/roundingadder/add_57/carry [3]) );
  XOR2X1 U7416 ( .IN1(
        \add_1_root_fmul_0_0_0_0_1/roundingadder/add_57/carry [2]), .IN2(
        \fmul_0_0_0_0_1/roundingadder/x_1_d1 [2]), .Q(\U503/DATA2_2 ) );
  AND2X1 U7417 ( .IN1(\fmul_0_0_0_0_1/roundingadder/x_1_d1 [1]), .IN2(
        \add_1_root_fmul_0_0_0_0_1/roundingadder/add_57/carry [1]), .Q(
        \add_1_root_fmul_0_0_0_0_1/roundingadder/add_57/carry [2]) );
  XOR2X1 U7418 ( .IN1(
        \add_1_root_fmul_0_0_0_0_1/roundingadder/add_57/carry [1]), .IN2(
        \fmul_0_0_0_0_1/roundingadder/x_1_d1 [1]), .Q(\U503/DATA2_1 ) );
  AND2X1 U7419 ( .IN1(\fmul_0_0_0_0_1/roundingadder/x_1_d1 [0]), .IN2(
        \fmul_0_0_0_0_1/roundingadder/n151_o[0] ), .Q(
        \add_1_root_fmul_0_0_0_0_1/roundingadder/add_57/carry [1]) );
  XOR2X1 U7420 ( .IN1(\fmul_0_0_0_0_1/roundingadder/n151_o[0] ), .IN2(
        \fmul_0_0_0_0_1/roundingadder/x_1_d1 [0]), .Q(\U503/DATA2_0 ) );
  XNOR2X1 U7421 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/A[5] ), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/carry [5]), .Q(
        \fmul_0_0_0_0_1/exppostnorm [5]) );
  OR2X1 U7422 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/carry [4]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/A[4] ), .Q(
        \add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/carry [5]) );
  XNOR2X1 U7423 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/A[4] ), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/carry [4]), .Q(
        \fmul_0_0_0_0_1/exppostnorm [4]) );
  AND2X1 U7424 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/carry [3]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/A[3] ), .Q(
        \add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/carry [4]) );
  XOR2X1 U7425 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/carry [3]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/A[3] ), .Q(
        \fmul_0_0_0_0_1/exppostnorm [3]) );
  AND2X1 U7426 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/carry [2]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/A[2] ), .Q(
        \add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/carry [3]) );
  XOR2X1 U7427 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/carry [2]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/A[2] ), .Q(
        \fmul_0_0_0_0_1/exppostnorm [2]) );
  AND2X1 U7428 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/B[0] ), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/A[0] ), .Q(
        \add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/carry [1]) );
  XOR2X1 U7429 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/B[0] ), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/A[0] ), .Q(
        \fmul_0_0_0_0_1/exppostnorm [0]) );
  AND2X1 U7430 ( .IN1(n5886), .IN2(n5874), .Q(
        \add_2_root_sub_1_root_fmul_0_0_0_0_1/add_321/carry [1]) );
  XOR2X1 U7431 ( .IN1(n5874), .IN2(n5886), .Q(
        \add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/A[0] ) );
  XNOR2X1 U7432 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/A[5] ), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/carry [5]), .Q(
        \fmul_0_0_0_0_0/exppostnorm [5]) );
  OR2X1 U7433 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/carry [4]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/A[4] ), .Q(
        \add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/carry [5]) );
  XNOR2X1 U7434 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/A[4] ), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/carry [4]), .Q(
        \fmul_0_0_0_0_0/exppostnorm [4]) );
  AND2X1 U7435 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/carry [3]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/A[3] ), .Q(
        \add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/carry [4]) );
  XOR2X1 U7436 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/carry [3]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/A[3] ), .Q(
        \fmul_0_0_0_0_0/exppostnorm [3]) );
  AND2X1 U7437 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/carry [2]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/A[2] ), .Q(
        \add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/carry [3]) );
  XOR2X1 U7438 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/carry [2]), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/A[2] ), .Q(
        \fmul_0_0_0_0_0/exppostnorm [2]) );
  AND2X1 U7439 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/B[0] ), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/A[0] ), .Q(
        \add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/carry [1]) );
  XOR2X1 U7440 ( .IN1(\add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/B[0] ), 
        .IN2(\add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/A[0] ), .Q(
        \fmul_0_0_0_0_0/exppostnorm [0]) );
  AND2X1 U7441 ( .IN1(n5958), .IN2(n5946), .Q(
        \add_2_root_sub_1_root_fmul_0_0_0_0_0/add_321/carry [1]) );
  XOR2X1 U7442 ( .IN1(n5946), .IN2(n5958), .Q(
        \add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/A[0] ) );
  AND2X1 U7443 ( .IN1(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[4] ), .IN2(n14516), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[5] ) );
  XOR2X1 U7444 ( .IN1(n14516), .IN2(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[4] ), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[4] ) );
  AND2X1 U7445 ( .IN1(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[3] ), .IN2(n14515), .Q(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[4] ) );
  XOR2X1 U7446 ( .IN1(n14515), .IN2(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[3] ), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[3] ) );
  AND2X1 U7447 ( .IN1(n14513), .IN2(n14514), .Q(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[3] ) );
  XOR2X1 U7448 ( .IN1(n14514), .IN2(n14513), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[2] ) );
  AND2X1 U7449 ( .IN1(
        \add_0_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .IN2(\fadd_0_0_0_0_9/fracyclose1 [1]), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [2]) );
  XOR2X1 U7450 ( .IN1(
        \add_0_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .IN2(\fadd_0_0_0_0_9/fracyclose1 [1]), .Q(\fadd_0_0_0_0_9/fracrcloseymx [1])
         );
  XNOR2X1 U7451 ( .IN1(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_9/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [5]), .IN2(n10654), .Q(\fadd_0_0_0_0_9/fracrclosexmy [5]) );
  OR2X1 U7452 ( .IN1(n14634), .IN2(n5346), .Q(
        \fadd_0_0_0_0_9/sub_707/carry [1]) );
  XNOR2X1 U7453 ( .IN1(n5346), .IN2(n14634), .Q(
        \fadd_0_0_0_0_9/exponentdifferencexy [0]) );
  OR2X1 U7454 ( .IN1(n14639), .IN2(n5334), .Q(
        \fadd_0_0_0_0_9/sub_710/carry [1]) );
  XNOR2X1 U7455 ( .IN1(n5334), .IN2(n14639), .Q(
        \fadd_0_0_0_0_9/exponentdifferenceyx [0]) );
  AND2X1 U7456 ( .IN1(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[4] ), .IN2(n14525), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[5] ) );
  XOR2X1 U7457 ( .IN1(n14525), .IN2(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[4] ), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[4] ) );
  AND2X1 U7458 ( .IN1(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[3] ), .IN2(n14524), .Q(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[4] ) );
  XOR2X1 U7459 ( .IN1(n14524), .IN2(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[3] ), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[3] ) );
  AND2X1 U7460 ( .IN1(n14522), .IN2(n14523), .Q(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[3] ) );
  XOR2X1 U7461 ( .IN1(n14523), .IN2(n14522), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[2] ) );
  AND2X1 U7462 ( .IN1(
        \add_0_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .IN2(\fadd_0_0_0_0_8/fracyclose1 [1]), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [2]) );
  XOR2X1 U7463 ( .IN1(
        \add_0_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .IN2(\fadd_0_0_0_0_8/fracyclose1 [1]), .Q(\fadd_0_0_0_0_8/fracrcloseymx [1])
         );
  XNOR2X1 U7464 ( .IN1(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_8/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [5]), .IN2(n10737), .Q(\fadd_0_0_0_0_8/fracrclosexmy [5]) );
  OR2X1 U7465 ( .IN1(n14623), .IN2(n5418), .Q(
        \fadd_0_0_0_0_8/sub_707/carry [1]) );
  XNOR2X1 U7466 ( .IN1(n5418), .IN2(n14623), .Q(
        \fadd_0_0_0_0_8/exponentdifferencexy [0]) );
  OR2X1 U7467 ( .IN1(n14628), .IN2(n5406), .Q(
        \fadd_0_0_0_0_8/sub_710/carry [1]) );
  XNOR2X1 U7468 ( .IN1(n5406), .IN2(n14628), .Q(
        \fadd_0_0_0_0_8/exponentdifferenceyx [0]) );
  AND2X1 U7469 ( .IN1(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[4] ), .IN2(n14480), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[5] ) );
  XOR2X1 U7470 ( .IN1(n14480), .IN2(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[4] ), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[4] ) );
  AND2X1 U7471 ( .IN1(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[3] ), .IN2(n14479), .Q(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[4] ) );
  XOR2X1 U7472 ( .IN1(n14479), .IN2(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[3] ), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[3] ) );
  AND2X1 U7473 ( .IN1(n14477), .IN2(n14478), .Q(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[3] ) );
  XOR2X1 U7474 ( .IN1(n14478), .IN2(n14477), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[2] ) );
  AND2X1 U7475 ( .IN1(
        \add_0_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .IN2(\fadd_0_0_0_0_7/fracyclose1 [1]), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [2]) );
  XOR2X1 U7476 ( .IN1(
        \add_0_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .IN2(\fadd_0_0_0_0_7/fracyclose1 [1]), .Q(\fadd_0_0_0_0_7/fracrcloseymx [1])
         );
  XNOR2X1 U7477 ( .IN1(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_7/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [5]), .IN2(n10818), .Q(\fadd_0_0_0_0_7/fracrclosexmy [5]) );
  OR2X1 U7478 ( .IN1(n14612), .IN2(n5490), .Q(
        \fadd_0_0_0_0_7/sub_707/carry [1]) );
  XNOR2X1 U7479 ( .IN1(n5490), .IN2(n14612), .Q(
        \fadd_0_0_0_0_7/exponentdifferencexy [0]) );
  OR2X1 U7480 ( .IN1(n14617), .IN2(n5478), .Q(
        \fadd_0_0_0_0_7/sub_710/carry [1]) );
  XNOR2X1 U7481 ( .IN1(n5478), .IN2(n14617), .Q(
        \fadd_0_0_0_0_7/exponentdifferenceyx [0]) );
  AND2X1 U7482 ( .IN1(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[4] ), .IN2(n14489), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[5] ) );
  XOR2X1 U7483 ( .IN1(n14489), .IN2(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[4] ), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[4] ) );
  AND2X1 U7484 ( .IN1(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[3] ), .IN2(n14488), .Q(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[4] ) );
  XOR2X1 U7485 ( .IN1(n14488), .IN2(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[3] ), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[3] ) );
  AND2X1 U7486 ( .IN1(n14486), .IN2(n14487), .Q(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[3] ) );
  XOR2X1 U7487 ( .IN1(n14487), .IN2(n14486), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[2] ) );
  AND2X1 U7488 ( .IN1(
        \add_0_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .IN2(\fadd_0_0_0_0_6/fracyclose1 [1]), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [2]) );
  XOR2X1 U7489 ( .IN1(
        \add_0_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .IN2(\fadd_0_0_0_0_6/fracyclose1 [1]), .Q(\fadd_0_0_0_0_6/fracrcloseymx [1])
         );
  XNOR2X1 U7490 ( .IN1(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_6/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [5]), .IN2(n10899), .Q(\fadd_0_0_0_0_6/fracrclosexmy [5]) );
  OR2X1 U7491 ( .IN1(n14601), .IN2(n5562), .Q(
        \fadd_0_0_0_0_6/sub_707/carry [1]) );
  XNOR2X1 U7492 ( .IN1(n5562), .IN2(n14601), .Q(
        \fadd_0_0_0_0_6/exponentdifferencexy [0]) );
  OR2X1 U7493 ( .IN1(n14606), .IN2(n5550), .Q(
        \fadd_0_0_0_0_6/sub_710/carry [1]) );
  XNOR2X1 U7494 ( .IN1(n5550), .IN2(n14606), .Q(
        \fadd_0_0_0_0_6/exponentdifferenceyx [0]) );
  AND2X1 U7495 ( .IN1(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[4] ), .IN2(n14471), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[5] ) );
  XOR2X1 U7496 ( .IN1(n14471), .IN2(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[4] ), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[4] ) );
  AND2X1 U7497 ( .IN1(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[3] ), .IN2(n14470), .Q(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[4] ) );
  XOR2X1 U7498 ( .IN1(n14470), .IN2(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[3] ), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[3] ) );
  AND2X1 U7499 ( .IN1(n14468), .IN2(n14469), .Q(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[3] ) );
  XOR2X1 U7500 ( .IN1(n14469), .IN2(n14468), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[2] ) );
  AND2X1 U7501 ( .IN1(
        \add_0_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .IN2(\fadd_0_0_0_0_5/fracyclose1 [1]), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [2]) );
  XOR2X1 U7502 ( .IN1(
        \add_0_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .IN2(\fadd_0_0_0_0_5/fracyclose1 [1]), .Q(\fadd_0_0_0_0_5/fracrcloseymx [1])
         );
  XNOR2X1 U7503 ( .IN1(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_5/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [5]), .IN2(n10980), .Q(\fadd_0_0_0_0_5/fracrclosexmy [5]) );
  OR2X1 U7504 ( .IN1(n14590), .IN2(n5634), .Q(
        \fadd_0_0_0_0_5/sub_707/carry [1]) );
  XNOR2X1 U7505 ( .IN1(n5634), .IN2(n14590), .Q(
        \fadd_0_0_0_0_5/exponentdifferencexy [0]) );
  OR2X1 U7506 ( .IN1(n14595), .IN2(n5622), .Q(
        \fadd_0_0_0_0_5/sub_710/carry [1]) );
  XNOR2X1 U7507 ( .IN1(n5622), .IN2(n14595), .Q(
        \fadd_0_0_0_0_5/exponentdifferenceyx [0]) );
  AND2X1 U7508 ( .IN1(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[4] ), .IN2(n14498), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[5] ) );
  XOR2X1 U7509 ( .IN1(n14498), .IN2(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[4] ), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[4] ) );
  AND2X1 U7510 ( .IN1(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[3] ), .IN2(n14497), .Q(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[4] ) );
  XOR2X1 U7511 ( .IN1(n14497), .IN2(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[3] ), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[3] ) );
  AND2X1 U7512 ( .IN1(n14495), .IN2(n14496), .Q(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[3] ) );
  XOR2X1 U7513 ( .IN1(n14496), .IN2(n14495), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[2] ) );
  AND2X1 U7514 ( .IN1(
        \add_0_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .IN2(\fadd_0_0_0_0_4/fracyclose1 [1]), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [2]) );
  XOR2X1 U7515 ( .IN1(
        \add_0_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .IN2(\fadd_0_0_0_0_4/fracyclose1 [1]), .Q(\fadd_0_0_0_0_4/fracrcloseymx [1])
         );
  XNOR2X1 U7516 ( .IN1(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_4/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [5]), .IN2(n11061), .Q(\fadd_0_0_0_0_4/fracrclosexmy [5]) );
  OR2X1 U7517 ( .IN1(n14579), .IN2(n5706), .Q(
        \fadd_0_0_0_0_4/sub_707/carry [1]) );
  XNOR2X1 U7518 ( .IN1(n5706), .IN2(n14579), .Q(
        \fadd_0_0_0_0_4/exponentdifferencexy [0]) );
  OR2X1 U7519 ( .IN1(n14584), .IN2(n5694), .Q(
        \fadd_0_0_0_0_4/sub_710/carry [1]) );
  XNOR2X1 U7520 ( .IN1(n5694), .IN2(n14584), .Q(
        \fadd_0_0_0_0_4/exponentdifferenceyx [0]) );
  AND2X1 U7521 ( .IN1(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[4] ), .IN2(n14453), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[5] ) );
  XOR2X1 U7522 ( .IN1(n14453), .IN2(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[4] ), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[4] ) );
  AND2X1 U7523 ( .IN1(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[3] ), .IN2(n14452), .Q(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[4] ) );
  XOR2X1 U7524 ( .IN1(n14452), .IN2(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[3] ), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[3] ) );
  AND2X1 U7525 ( .IN1(n14450), .IN2(n14451), .Q(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[3] ) );
  XOR2X1 U7526 ( .IN1(n14451), .IN2(n14450), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[2] ) );
  AND2X1 U7527 ( .IN1(
        \add_0_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .IN2(\fadd_0_0_0_0_3/fracyclose1 [1]), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [2]) );
  XOR2X1 U7528 ( .IN1(
        \add_0_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .IN2(\fadd_0_0_0_0_3/fracyclose1 [1]), .Q(\fadd_0_0_0_0_3/fracrcloseymx [1])
         );
  XNOR2X1 U7529 ( .IN1(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_3/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [5]), .IN2(n11142), .Q(\fadd_0_0_0_0_3/fracrclosexmy [5]) );
  OR2X1 U7530 ( .IN1(n14568), .IN2(n5778), .Q(
        \fadd_0_0_0_0_3/sub_707/carry [1]) );
  XNOR2X1 U7531 ( .IN1(n5778), .IN2(n14568), .Q(
        \fadd_0_0_0_0_3/exponentdifferencexy [0]) );
  OR2X1 U7532 ( .IN1(n14573), .IN2(n5766), .Q(
        \fadd_0_0_0_0_3/sub_710/carry [1]) );
  XNOR2X1 U7533 ( .IN1(n5766), .IN2(n14573), .Q(
        \fadd_0_0_0_0_3/exponentdifferenceyx [0]) );
  AND2X1 U7534 ( .IN1(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[4] ), .IN2(n14462), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[5] ) );
  XOR2X1 U7535 ( .IN1(n14462), .IN2(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[4] ), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[4] ) );
  AND2X1 U7536 ( .IN1(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[3] ), .IN2(n14461), .Q(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[4] ) );
  XOR2X1 U7537 ( .IN1(n14461), .IN2(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[3] ), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[3] ) );
  AND2X1 U7538 ( .IN1(n14459), .IN2(n14460), .Q(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[3] ) );
  XOR2X1 U7539 ( .IN1(n14460), .IN2(n14459), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[2] ) );
  AND2X1 U7540 ( .IN1(
        \add_0_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .IN2(\fadd_0_0_0_0_2/fracyclose1 [1]), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [2]) );
  XOR2X1 U7541 ( .IN1(
        \add_0_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .IN2(\fadd_0_0_0_0_2/fracyclose1 [1]), .Q(\fadd_0_0_0_0_2/fracrcloseymx [1])
         );
  XNOR2X1 U7542 ( .IN1(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_2/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [5]), .IN2(n11223), .Q(\fadd_0_0_0_0_2/fracrclosexmy [5]) );
  OR2X1 U7543 ( .IN1(n14557), .IN2(n5850), .Q(
        \fadd_0_0_0_0_2/sub_707/carry [1]) );
  XNOR2X1 U7544 ( .IN1(n5850), .IN2(n14557), .Q(
        \fadd_0_0_0_0_2/exponentdifferencexy [0]) );
  OR2X1 U7545 ( .IN1(n14561), .IN2(n5838), .Q(
        \fadd_0_0_0_0_2/sub_710/carry [1]) );
  XNOR2X1 U7546 ( .IN1(n5838), .IN2(n14561), .Q(
        \fadd_0_0_0_0_2/exponentdifferenceyx [0]) );
  AND2X1 U7547 ( .IN1(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[4] ), .IN2(n14444), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[5] ) );
  XOR2X1 U7548 ( .IN1(n14444), .IN2(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[4] ), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[4] ) );
  AND2X1 U7549 ( .IN1(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[3] ), .IN2(n14443), .Q(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[4] ) );
  XOR2X1 U7550 ( .IN1(n14443), .IN2(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[3] ), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[3] ) );
  AND2X1 U7551 ( .IN1(n14441), .IN2(n14442), .Q(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[3] ) );
  XOR2X1 U7552 ( .IN1(n14442), .IN2(n14441), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[2] ) );
  AND2X1 U7553 ( .IN1(
        \add_0_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .IN2(\fadd_0_0_0_0_1/fracyclose1 [1]), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [2]) );
  XOR2X1 U7554 ( .IN1(
        \add_0_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .IN2(\fadd_0_0_0_0_1/fracyclose1 [1]), .Q(\fadd_0_0_0_0_1/fracrcloseymx [1])
         );
  XNOR2X1 U7555 ( .IN1(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_1/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [5]), .IN2(n11359), .Q(\fadd_0_0_0_0_1/fracrclosexmy [5]) );
  OR2X1 U7556 ( .IN1(n14546), .IN2(n5922), .Q(
        \fadd_0_0_0_0_1/sub_707/carry [1]) );
  XNOR2X1 U7557 ( .IN1(n5922), .IN2(n14546), .Q(
        \fadd_0_0_0_0_1/exponentdifferencexy [0]) );
  OR2X1 U7558 ( .IN1(n14551), .IN2(n5910), .Q(
        \fadd_0_0_0_0_1/sub_710/carry [1]) );
  XNOR2X1 U7559 ( .IN1(n5910), .IN2(n14551), .Q(
        \fadd_0_0_0_0_1/exponentdifferenceyx [0]) );
  AND2X1 U7560 ( .IN1(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[4] ), .IN2(n14507), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[5] ) );
  XOR2X1 U7561 ( .IN1(n14507), .IN2(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[4] ), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[4] ) );
  AND2X1 U7562 ( .IN1(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[3] ), .IN2(n14506), .Q(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[4] ) );
  XOR2X1 U7563 ( .IN1(n14506), .IN2(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[3] ), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[3] ) );
  AND2X1 U7564 ( .IN1(n14504), .IN2(n14505), .Q(
        \sub_2_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry[3] ) );
  XOR2X1 U7565 ( .IN1(n14505), .IN2(n14504), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[2] ) );
  AND2X1 U7566 ( .IN1(
        \add_0_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .IN2(\fadd_0_0_0_0_0/fracyclose1 [1]), .Q(
        \add_0_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_303/carry [2]) );
  XOR2X1 U7567 ( .IN1(
        \add_0_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_303/B[1] ), .IN2(\fadd_0_0_0_0_0/fracyclose1 [1]), .Q(\fadd_0_0_0_0_0/fracrcloseymx [1])
         );
  XNOR2X1 U7568 ( .IN1(
        \sub_0_root_sub_1_root_fadd_0_0_0_0_0/fpadd_5_4_f300_uid2_dualsubclose/add_300/carry [5]), .IN2(n11442), .Q(\fadd_0_0_0_0_0/fracrclosexmy [5]) );
  OR2X1 U7569 ( .IN1(n14535), .IN2(n5994), .Q(
        \fadd_0_0_0_0_0/sub_707/carry [1]) );
  XNOR2X1 U7570 ( .IN1(n5994), .IN2(n14535), .Q(
        \fadd_0_0_0_0_0/exponentdifferencexy [0]) );
  OR2X1 U7571 ( .IN1(n14540), .IN2(n5982), .Q(
        \fadd_0_0_0_0_0/sub_710/carry [1]) );
  XNOR2X1 U7572 ( .IN1(n5982), .IN2(n14540), .Q(
        \fadd_0_0_0_0_0/exponentdifferenceyx [0]) );
  INVX0 U7573 ( .INP(\add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/B[1] ), 
        .ZN(\add_0_root_sub_1_root_fmul_0_0_0_0_9/add_321/B[0] ) );
  INVX0 U7574 ( .INP(\add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/B[1] ), 
        .ZN(\add_0_root_sub_1_root_fmul_0_0_0_0_8/add_321/B[0] ) );
  INVX0 U7575 ( .INP(\add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/B[1] ), 
        .ZN(\add_0_root_sub_1_root_fmul_0_0_0_0_7/add_321/B[0] ) );
  INVX0 U7576 ( .INP(\add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/B[1] ), 
        .ZN(\add_0_root_sub_1_root_fmul_0_0_0_0_6/add_321/B[0] ) );
  INVX0 U7577 ( .INP(\add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/B[1] ), 
        .ZN(\add_0_root_sub_1_root_fmul_0_0_0_0_5/add_321/B[0] ) );
  INVX0 U7578 ( .INP(\add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/B[1] ), 
        .ZN(\add_0_root_sub_1_root_fmul_0_0_0_0_4/add_321/B[0] ) );
  INVX0 U7579 ( .INP(\add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/B[1] ), 
        .ZN(\add_0_root_sub_1_root_fmul_0_0_0_0_3/add_321/B[0] ) );
  INVX0 U7580 ( .INP(\add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/B[1] ), 
        .ZN(\add_0_root_sub_1_root_fmul_0_0_0_0_2/add_321/B[0] ) );
  INVX0 U7581 ( .INP(\add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/B[1] ), 
        .ZN(\add_0_root_sub_1_root_fmul_0_0_0_0_1/add_321/B[0] ) );
  INVX0 U7582 ( .INP(\add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/B[1] ), 
        .ZN(\add_0_root_sub_1_root_fmul_0_0_0_0_0/add_321/B[0] ) );
  INVX0 U7583 ( .INP(\fadd_0_0_0_0_0/sub_707/carry [5]), .ZN(
        \fadd_0_0_0_0_0/exponentdifferencexy [5]) );
  INVX0 U7584 ( .INP(\fadd_0_0_0_0_1/sub_707/carry [5]), .ZN(
        \fadd_0_0_0_0_1/exponentdifferencexy [5]) );
  INVX0 U7585 ( .INP(\fadd_0_0_0_0_2/sub_707/carry [5]), .ZN(
        \fadd_0_0_0_0_2/exponentdifferencexy [5]) );
  INVX0 U7586 ( .INP(\fadd_0_0_0_0_3/sub_707/carry [5]), .ZN(
        \fadd_0_0_0_0_3/exponentdifferencexy [5]) );
  INVX0 U7587 ( .INP(\fadd_0_0_0_0_4/sub_707/carry [5]), .ZN(
        \fadd_0_0_0_0_4/exponentdifferencexy [5]) );
  INVX0 U7588 ( .INP(\fadd_0_0_0_0_5/sub_707/carry [5]), .ZN(
        \fadd_0_0_0_0_5/exponentdifferencexy [5]) );
  INVX0 U7589 ( .INP(\fadd_0_0_0_0_6/sub_707/carry [5]), .ZN(
        \fadd_0_0_0_0_6/exponentdifferencexy [5]) );
  INVX0 U7590 ( .INP(\fadd_0_0_0_0_7/sub_707/carry [5]), .ZN(
        \fadd_0_0_0_0_7/exponentdifferencexy [5]) );
  INVX0 U7591 ( .INP(\fadd_0_0_0_0_8/sub_707/carry [5]), .ZN(
        \fadd_0_0_0_0_8/exponentdifferencexy [5]) );
  INVX0 U7592 ( .INP(\fadd_0_0_0_0_9/sub_707/carry [5]), .ZN(
        \fadd_0_0_0_0_9/exponentdifferencexy [5]) );
endmodule

