`default_nettype none
module linear (
	clk,
	rst,
	p__arg0_0_0,
	p__arg0_0_1,
	p__arg0_0_10,
	p__arg0_0_2,
	p__arg0_0_3,
	p__arg0_0_4,
	p__arg0_0_5,
	p__arg0_0_6,
	p__arg0_0_7,
	p__arg0_0_8,
	p__arg0_0_9,
	p___constant_11x11xf32_0_0,
	p___constant_11x11xf32_0_1,
	p___constant_11x11xf32_0_10,
	p___constant_11x11xf32_0_2,
	p___constant_11x11xf32_0_3,
	p___constant_11x11xf32_0_4,
	p___constant_11x11xf32_0_5,
	p___constant_11x11xf32_0_6,
	p___constant_11x11xf32_0_7,
	p___constant_11x11xf32_0_8,
	p___constant_11x11xf32_0_9,
	p___constant_11x11xf32_10_0,
	p___constant_11x11xf32_10_1,
	p___constant_11x11xf32_10_10,
	p___constant_11x11xf32_10_2,
	p___constant_11x11xf32_10_3,
	p___constant_11x11xf32_10_4,
	p___constant_11x11xf32_10_5,
	p___constant_11x11xf32_10_6,
	p___constant_11x11xf32_10_7,
	p___constant_11x11xf32_10_8,
	p___constant_11x11xf32_10_9,
	p___constant_11x11xf32_1_0,
	p___constant_11x11xf32_1_1,
	p___constant_11x11xf32_1_10,
	p___constant_11x11xf32_1_2,
	p___constant_11x11xf32_1_3,
	p___constant_11x11xf32_1_4,
	p___constant_11x11xf32_1_5,
	p___constant_11x11xf32_1_6,
	p___constant_11x11xf32_1_7,
	p___constant_11x11xf32_1_8,
	p___constant_11x11xf32_1_9,
	p___constant_11x11xf32_2_0,
	p___constant_11x11xf32_2_1,
	p___constant_11x11xf32_2_10,
	p___constant_11x11xf32_2_2,
	p___constant_11x11xf32_2_3,
	p___constant_11x11xf32_2_4,
	p___constant_11x11xf32_2_5,
	p___constant_11x11xf32_2_6,
	p___constant_11x11xf32_2_7,
	p___constant_11x11xf32_2_8,
	p___constant_11x11xf32_2_9,
	p___constant_11x11xf32_3_0,
	p___constant_11x11xf32_3_1,
	p___constant_11x11xf32_3_10,
	p___constant_11x11xf32_3_2,
	p___constant_11x11xf32_3_3,
	p___constant_11x11xf32_3_4,
	p___constant_11x11xf32_3_5,
	p___constant_11x11xf32_3_6,
	p___constant_11x11xf32_3_7,
	p___constant_11x11xf32_3_8,
	p___constant_11x11xf32_3_9,
	p___constant_11x11xf32_4_0,
	p___constant_11x11xf32_4_1,
	p___constant_11x11xf32_4_10,
	p___constant_11x11xf32_4_2,
	p___constant_11x11xf32_4_3,
	p___constant_11x11xf32_4_4,
	p___constant_11x11xf32_4_5,
	p___constant_11x11xf32_4_6,
	p___constant_11x11xf32_4_7,
	p___constant_11x11xf32_4_8,
	p___constant_11x11xf32_4_9,
	p___constant_11x11xf32_5_0,
	p___constant_11x11xf32_5_1,
	p___constant_11x11xf32_5_10,
	p___constant_11x11xf32_5_2,
	p___constant_11x11xf32_5_3,
	p___constant_11x11xf32_5_4,
	p___constant_11x11xf32_5_5,
	p___constant_11x11xf32_5_6,
	p___constant_11x11xf32_5_7,
	p___constant_11x11xf32_5_8,
	p___constant_11x11xf32_5_9,
	p___constant_11x11xf32_6_0,
	p___constant_11x11xf32_6_1,
	p___constant_11x11xf32_6_10,
	p___constant_11x11xf32_6_2,
	p___constant_11x11xf32_6_3,
	p___constant_11x11xf32_6_4,
	p___constant_11x11xf32_6_5,
	p___constant_11x11xf32_6_6,
	p___constant_11x11xf32_6_7,
	p___constant_11x11xf32_6_8,
	p___constant_11x11xf32_6_9,
	p___constant_11x11xf32_7_0,
	p___constant_11x11xf32_7_1,
	p___constant_11x11xf32_7_10,
	p___constant_11x11xf32_7_2,
	p___constant_11x11xf32_7_3,
	p___constant_11x11xf32_7_4,
	p___constant_11x11xf32_7_5,
	p___constant_11x11xf32_7_6,
	p___constant_11x11xf32_7_7,
	p___constant_11x11xf32_7_8,
	p___constant_11x11xf32_7_9,
	p___constant_11x11xf32_8_0,
	p___constant_11x11xf32_8_1,
	p___constant_11x11xf32_8_10,
	p___constant_11x11xf32_8_2,
	p___constant_11x11xf32_8_3,
	p___constant_11x11xf32_8_4,
	p___constant_11x11xf32_8_5,
	p___constant_11x11xf32_8_6,
	p___constant_11x11xf32_8_7,
	p___constant_11x11xf32_8_8,
	p___constant_11x11xf32_8_9,
	p___constant_11x11xf32_9_0,
	p___constant_11x11xf32_9_1,
	p___constant_11x11xf32_9_10,
	p___constant_11x11xf32_9_2,
	p___constant_11x11xf32_9_3,
	p___constant_11x11xf32_9_4,
	p___constant_11x11xf32_9_5,
	p___constant_11x11xf32_9_6,
	p___constant_11x11xf32_9_7,
	p___constant_11x11xf32_9_8,
	p___constant_11x11xf32_9_9,
	p___constant_11xf32_0,
	p___constant_11xf32_1,
	p___constant_11xf32_10,
	p___constant_11xf32_2,
	p___constant_11xf32_3,
	p___constant_11xf32_4,
	p___constant_11xf32_5,
	p___constant_11xf32_6,
	p___constant_11xf32_7,
	p___constant_11xf32_8,
	p___constant_11xf32_9,
	output_p_val_313
);
	input wire clk;
	input wire rst;
	input wire [11:0] p__arg0_0_0;
	input wire [11:0] p__arg0_0_1;
	input wire [11:0] p__arg0_0_10;
	input wire [11:0] p__arg0_0_2;
	input wire [11:0] p__arg0_0_3;
	input wire [11:0] p__arg0_0_4;
	input wire [11:0] p__arg0_0_5;
	input wire [11:0] p__arg0_0_6;
	input wire [11:0] p__arg0_0_7;
	input wire [11:0] p__arg0_0_8;
	input wire [11:0] p__arg0_0_9;
	input wire [11:0] p___constant_11x11xf32_0_0;
	input wire [11:0] p___constant_11x11xf32_0_1;
	input wire [11:0] p___constant_11x11xf32_0_10;
	input wire [11:0] p___constant_11x11xf32_0_2;
	input wire [11:0] p___constant_11x11xf32_0_3;
	input wire [11:0] p___constant_11x11xf32_0_4;
	input wire [11:0] p___constant_11x11xf32_0_5;
	input wire [11:0] p___constant_11x11xf32_0_6;
	input wire [11:0] p___constant_11x11xf32_0_7;
	input wire [11:0] p___constant_11x11xf32_0_8;
	input wire [11:0] p___constant_11x11xf32_0_9;
	input wire [11:0] p___constant_11x11xf32_10_0;
	input wire [11:0] p___constant_11x11xf32_10_1;
	input wire [11:0] p___constant_11x11xf32_10_10;
	input wire [11:0] p___constant_11x11xf32_10_2;
	input wire [11:0] p___constant_11x11xf32_10_3;
	input wire [11:0] p___constant_11x11xf32_10_4;
	input wire [11:0] p___constant_11x11xf32_10_5;
	input wire [11:0] p___constant_11x11xf32_10_6;
	input wire [11:0] p___constant_11x11xf32_10_7;
	input wire [11:0] p___constant_11x11xf32_10_8;
	input wire [11:0] p___constant_11x11xf32_10_9;
	input wire [11:0] p___constant_11x11xf32_1_0;
	input wire [11:0] p___constant_11x11xf32_1_1;
	input wire [11:0] p___constant_11x11xf32_1_10;
	input wire [11:0] p___constant_11x11xf32_1_2;
	input wire [11:0] p___constant_11x11xf32_1_3;
	input wire [11:0] p___constant_11x11xf32_1_4;
	input wire [11:0] p___constant_11x11xf32_1_5;
	input wire [11:0] p___constant_11x11xf32_1_6;
	input wire [11:0] p___constant_11x11xf32_1_7;
	input wire [11:0] p___constant_11x11xf32_1_8;
	input wire [11:0] p___constant_11x11xf32_1_9;
	input wire [11:0] p___constant_11x11xf32_2_0;
	input wire [11:0] p___constant_11x11xf32_2_1;
	input wire [11:0] p___constant_11x11xf32_2_10;
	input wire [11:0] p___constant_11x11xf32_2_2;
	input wire [11:0] p___constant_11x11xf32_2_3;
	input wire [11:0] p___constant_11x11xf32_2_4;
	input wire [11:0] p___constant_11x11xf32_2_5;
	input wire [11:0] p___constant_11x11xf32_2_6;
	input wire [11:0] p___constant_11x11xf32_2_7;
	input wire [11:0] p___constant_11x11xf32_2_8;
	input wire [11:0] p___constant_11x11xf32_2_9;
	input wire [11:0] p___constant_11x11xf32_3_0;
	input wire [11:0] p___constant_11x11xf32_3_1;
	input wire [11:0] p___constant_11x11xf32_3_10;
	input wire [11:0] p___constant_11x11xf32_3_2;
	input wire [11:0] p___constant_11x11xf32_3_3;
	input wire [11:0] p___constant_11x11xf32_3_4;
	input wire [11:0] p___constant_11x11xf32_3_5;
	input wire [11:0] p___constant_11x11xf32_3_6;
	input wire [11:0] p___constant_11x11xf32_3_7;
	input wire [11:0] p___constant_11x11xf32_3_8;
	input wire [11:0] p___constant_11x11xf32_3_9;
	input wire [11:0] p___constant_11x11xf32_4_0;
	input wire [11:0] p___constant_11x11xf32_4_1;
	input wire [11:0] p___constant_11x11xf32_4_10;
	input wire [11:0] p___constant_11x11xf32_4_2;
	input wire [11:0] p___constant_11x11xf32_4_3;
	input wire [11:0] p___constant_11x11xf32_4_4;
	input wire [11:0] p___constant_11x11xf32_4_5;
	input wire [11:0] p___constant_11x11xf32_4_6;
	input wire [11:0] p___constant_11x11xf32_4_7;
	input wire [11:0] p___constant_11x11xf32_4_8;
	input wire [11:0] p___constant_11x11xf32_4_9;
	input wire [11:0] p___constant_11x11xf32_5_0;
	input wire [11:0] p___constant_11x11xf32_5_1;
	input wire [11:0] p___constant_11x11xf32_5_10;
	input wire [11:0] p___constant_11x11xf32_5_2;
	input wire [11:0] p___constant_11x11xf32_5_3;
	input wire [11:0] p___constant_11x11xf32_5_4;
	input wire [11:0] p___constant_11x11xf32_5_5;
	input wire [11:0] p___constant_11x11xf32_5_6;
	input wire [11:0] p___constant_11x11xf32_5_7;
	input wire [11:0] p___constant_11x11xf32_5_8;
	input wire [11:0] p___constant_11x11xf32_5_9;
	input wire [11:0] p___constant_11x11xf32_6_0;
	input wire [11:0] p___constant_11x11xf32_6_1;
	input wire [11:0] p___constant_11x11xf32_6_10;
	input wire [11:0] p___constant_11x11xf32_6_2;
	input wire [11:0] p___constant_11x11xf32_6_3;
	input wire [11:0] p___constant_11x11xf32_6_4;
	input wire [11:0] p___constant_11x11xf32_6_5;
	input wire [11:0] p___constant_11x11xf32_6_6;
	input wire [11:0] p___constant_11x11xf32_6_7;
	input wire [11:0] p___constant_11x11xf32_6_8;
	input wire [11:0] p___constant_11x11xf32_6_9;
	input wire [11:0] p___constant_11x11xf32_7_0;
	input wire [11:0] p___constant_11x11xf32_7_1;
	input wire [11:0] p___constant_11x11xf32_7_10;
	input wire [11:0] p___constant_11x11xf32_7_2;
	input wire [11:0] p___constant_11x11xf32_7_3;
	input wire [11:0] p___constant_11x11xf32_7_4;
	input wire [11:0] p___constant_11x11xf32_7_5;
	input wire [11:0] p___constant_11x11xf32_7_6;
	input wire [11:0] p___constant_11x11xf32_7_7;
	input wire [11:0] p___constant_11x11xf32_7_8;
	input wire [11:0] p___constant_11x11xf32_7_9;
	input wire [11:0] p___constant_11x11xf32_8_0;
	input wire [11:0] p___constant_11x11xf32_8_1;
	input wire [11:0] p___constant_11x11xf32_8_10;
	input wire [11:0] p___constant_11x11xf32_8_2;
	input wire [11:0] p___constant_11x11xf32_8_3;
	input wire [11:0] p___constant_11x11xf32_8_4;
	input wire [11:0] p___constant_11x11xf32_8_5;
	input wire [11:0] p___constant_11x11xf32_8_6;
	input wire [11:0] p___constant_11x11xf32_8_7;
	input wire [11:0] p___constant_11x11xf32_8_8;
	input wire [11:0] p___constant_11x11xf32_8_9;
	input wire [11:0] p___constant_11x11xf32_9_0;
	input wire [11:0] p___constant_11x11xf32_9_1;
	input wire [11:0] p___constant_11x11xf32_9_10;
	input wire [11:0] p___constant_11x11xf32_9_2;
	input wire [11:0] p___constant_11x11xf32_9_3;
	input wire [11:0] p___constant_11x11xf32_9_4;
	input wire [11:0] p___constant_11x11xf32_9_5;
	input wire [11:0] p___constant_11x11xf32_9_6;
	input wire [11:0] p___constant_11x11xf32_9_7;
	input wire [11:0] p___constant_11x11xf32_9_8;
	input wire [11:0] p___constant_11x11xf32_9_9;
	input wire [11:0] p___constant_11xf32_0;
	input wire [11:0] p___constant_11xf32_1;
	input wire [11:0] p___constant_11xf32_10;
	input wire [11:0] p___constant_11xf32_2;
	input wire [11:0] p___constant_11xf32_3;
	input wire [11:0] p___constant_11xf32_4;
	input wire [11:0] p___constant_11xf32_5;
	input wire [11:0] p___constant_11xf32_6;
	input wire [11:0] p___constant_11xf32_7;
	input wire [11:0] p___constant_11xf32_8;
	input wire [11:0] p___constant_11xf32_9;
	output wire [11:0] output_p_val_313;



endmodule

